library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_arith.all;

entity tb_axis_iic_bridge is 
end tb_axis_iic_bridge;



architecture tb_axis_iic_bridge_arch of tb_axis_iic_bridge is 

    constant N_BYTES            :           integer     := 4                                    ;
    constant CLK_PERIOD         :           integer     := 5000000                              ;
    constant CLK_I2C_PERIOD     :           integer     := 400000                               ; -- 4

    component axis_iic_ctrlr 
        generic (
            CLK_PERIOD      :           integer := 100000000                            ;
            CLK_I2C_PERIOD  :           integer := 400000                               ;
            N_BYTES         :           integer := 32                                   ;
            DEPTH           :           integer := 16                                    
        );  
        port (
            clk             :   in      std_logic                                       ;
            resetn          :   in      std_logic                                       ;
            s_axis_tdata    :   in      std_logic_vector ( ((N_BYTES*8)-1) downto 0 )   ;
            s_axis_tkeep    :   in      std_logic_vector (       N_BYTES-1 downto 0 )   ;
            s_axis_tdest    :   in      std_logic_vector (               7 downto 0 )   ;
            s_axis_tvalid   :   in      std_logic                                       ;
            s_axis_tready   :   out     std_logic                                       ;
            s_axis_tlast    :   in      std_logic                                       ;
            m_axis_tdata    :   out     std_logic_vector ( ((N_BYTES*8)-1) downto 0 )   ;
            m_axis_tkeep    :   out     std_logic_vector (       N_BYTES-1 downto 0 )   ;
            m_axis_tdest    :   out     std_logic_vector (               7 downto 0 )   ;
            m_axis_tvalid   :   out     std_logic                                       ;
            m_axis_tready   :   in      std_logic                                       ;
            m_axis_tlast    :   out     std_logic                                       ;
            scl_i           :   in      std_logic                                       ;
            sda_i           :   in      std_logic                                       ;
            scl_t           :   out     std_logic                                       ;
            sda_t           :   out     std_logic                                        
        );
    end component;

    component axis_iic_bridge 
        generic (
            CLK_PERIOD      :           integer     := 100000000                            ;
            CLK_I2C_PERIOD  :           integer     := 25000000                             ;
            N_BYTES         :           integer     := 32                                   ;
            WRITE_CONTROL   :           string      := "STREAM" -- or "COUNTER"
        ); 
        port (
            CLK             :   in      std_Logic                                           ;
            reset           :   in      std_Logic                                           ;
            s_axis_tdata    :   in      std_logic_Vector ( ((N_BYTES*8)-1) downto 0 )       ;
            s_axis_tkeep    :   in      std_logic_Vector (       N_BYTES-1 downto 0 )       ;
            s_axis_tuser    :   in      std_logic_Vector ( 7 downto 0 )                     ;
            s_axis_tvalid   :   in      std_Logic                                           ;
            s_axis_tready   :   out     std_Logic                                           ;
            s_axis_tlast    :   in      std_Logic                                           ;
            m_axis_tdata    :   out     std_logic_Vector ( ((N_BYTES*8)-1) downto 0 )       ;
            m_axis_tkeep    :   out     std_logic_Vector (       N_BYTES-1 downto 0 )       ;
            m_axis_tuser    :   out     std_logic_Vector ( 7 downto 0 )                     ;
            m_axis_tvalid   :   out     std_Logic                                           ;
            m_axis_tready   :   in      std_Logic                                           ;
            m_axis_tlast    :   out     std_Logic                                           ;
            scl_i           :   in      std_Logic                                           ;
            sda_i           :   in      std_Logic                                           ;
            scl_t           :   out     std_Logic                                           ;
            sda_t           :   out     std_Logic                                            
        );
    end component;


    signal  CLK             :           std_Logic                                     := '0'                ;
    signal  reset           :           std_Logic                                     := '0'                ;
    signal  s_axis_tdata    :           std_logic_Vector ( ((N_BYTES*8)-1) downto 0 ) := (others => '0')    ;
    signal  s_axis_tkeep    :           std_logic_Vector (       N_BYTES-1 downto 0 ) := (others => '0')    ;
    signal  s_axis_tuser    :           std_Logic_Vector (               7 downto 0 ) := (others => '0')    ;
    signal  s_axis_tvalid   :           std_Logic                                     := '0'                ;
    signal  s_axis_tready   :           std_Logic                                                           ;
    signal  s_axis_tlast    :           std_Logic                                     := '0'                ;

    signal  m_axis_tdata     :           std_logic_Vector ( ((N_BYTES*8)-1) downto 0 )                       ;
    signal  m_axis_tkeep     :           std_logic_Vector (       N_BYTES-1 downto 0 )                       ;
    signal  m_axis_tuser     :           std_Logic_Vector (               7 downto 0 )                       ;
    signal  m_axis_tvalid    :           std_Logic                                                           ;
    signal  m_axis_tready    :           std_Logic                                     := '0'                ;
    signal  m_axis_tlast     :           std_Logic                                                           ;


    signal  scl_i           :           std_Logic                                     := '0'                ;
    signal  sda_i           :           std_Logic                                     := '0'                ;
    signal  scl_t           :           std_Logic                                                           ;
    signal  sda_t           :           std_Logic                                                           ;

    constant clock_period   :           time                                          := 200 ns              ;

    signal i                :           integer                                       := 0                  ;

begin 

    CLK <= not CLK after clock_period/2;

    i_processing : process(CLK)
    begin
        if CLK'event AND CLK = '1' then 
            i <= i + 1;
        end if;
    end process;

    reset <= '1' when i < 5 else '0';

    s_axis_processing : process(CLK)
    begin
        if CLK'event AND CLK = '1' then 
            case i is
                when 100 => S_AXIS_TDATA <= x"00000039"; S_AXIS_TUSER <= x"A7"; S_AXIS_TKEEP <= "1111"; S_AXIS_TVALID <= '1'; S_AXIS_TLAST <= '1';
                when others => S_AXIS_TDATA <= S_AXIS_TDATA; S_AXIS_TUSER <= S_AXIS_TUSER; S_AXIS_TKEEP <= S_AXIS_TKEEP; S_AXIS_TVALID <= '0'; S_AXIS_TLAST <= S_AXIS_TLAST;
            end case;
        end if;
    end process;

    axis_iic_bridge_inst : axis_iic_bridge 
        generic map (
            CLK_PERIOD      =>  CLK_PERIOD                      ,
            CLK_I2C_PERIOD  =>  CLK_I2C_PERIOD                  ,
            N_BYTES         =>  N_BYTES                         ,
            WRITE_CONTROL   =>  "STREAM" -- or "COUNTER"
        )
        port map  (
            CLK             =>  CLK                             ,
            reset           =>  reset                           ,
            s_axis_tdata    =>  s_axis_tdata                    ,
            s_axis_tuser    =>  s_axis_tuser                    ,
            s_axis_tkeep    =>  s_axis_tkeep                    ,
            s_axis_tvalid   =>  s_axis_tvalid                   ,
            s_axis_tready   =>  open                            ,
            s_axis_tlast    =>  s_axis_tlast                    ,
            m_axis_tdata    =>  m_axis_tdata                    ,
            m_axis_tkeep    =>  m_axis_tkeep                    ,
            m_axis_tuser    =>  m_axis_tuser                    ,
            m_axis_tvalid   =>  m_axis_tvalid                   ,
            m_axis_tready   =>  m_axis_tready                   ,
            m_axis_tlast    =>  m_axis_tlast                    ,
            scl_i           =>  scl_i                           ,
            sda_i           =>  sda_i                           ,
            scl_t           =>  scl_t                           ,
            sda_t           =>  sda_t                            
        );

    scl_i <= scl_t;

    m_axis_tready <= '1';

    sda_i_processing : process(CLK)
    begin

        if CLK'event AND CLK = '1' then 
            case i is 
                when 0   => sda_i <= '1';

                when 107 => sda_i <= '1';
                when 108 => sda_i <= '0';
                when 109 => sda_i <= '0';
                when 110 => sda_i <= '0';
                when 111 => sda_i <= '0';
                when 112 => sda_i <= '0';
                when 113 => sda_i <= '0';
                when 114 => sda_i <= '0';
                when 115 => sda_i <= '0';
                when 116 => sda_i <= '0';
                when 117 => sda_i <= '0';
                when 118 => sda_i <= '0';
                when 119 => sda_i <= '0';
                when 120 => sda_i <= '1';
                when 121 => sda_i <= '1';
                when 122 => sda_i <= '1';
                when 123 => sda_i <= '1';
                when 124 => sda_i <= '1';
                when 125 => sda_i <= '1';
                when 126 => sda_i <= '1';
                when 127 => sda_i <= '1';
                when 128 => sda_i <= '1';
                when 129 => sda_i <= '1';
                when 130 => sda_i <= '1';
                when 131 => sda_i <= '1';
                when 132 => sda_i <= '0';
                when 133 => sda_i <= '0';
                when 134 => sda_i <= '0';
                when 135 => sda_i <= '0';
                when 136 => sda_i <= '0';
                when 137 => sda_i <= '0';
                when 138 => sda_i <= '0';
                when 139 => sda_i <= '0';
                when 140 => sda_i <= '0';
                when 141 => sda_i <= '0';
                when 142 => sda_i <= '0';
                when 143 => sda_i <= '0';
                when 144 => sda_i <= '1';
                when 145 => sda_i <= '1';
                when 146 => sda_i <= '1';
                when 147 => sda_i <= '1';
                when 148 => sda_i <= '1';
                when 149 => sda_i <= '1';
                when 150 => sda_i <= '1';
                when 151 => sda_i <= '1';
                when 152 => sda_i <= '1';
                when 153 => sda_i <= '1';
                when 154 => sda_i <= '1';
                when 155 => sda_i <= '1';
                when 156 => sda_i <= '0';
                when 157 => sda_i <= '0';
                when 158 => sda_i <= '0';
                when 159 => sda_i <= '0';
                when 160 => sda_i <= '0';
                when 161 => sda_i <= '0';
                when 162 => sda_i <= '0';
                when 163 => sda_i <= '0';
                when 164 => sda_i <= '0';
                when 165 => sda_i <= '0';
                when 166 => sda_i <= '0';
                when 167 => sda_i <= '0';
                when 168 => sda_i <= '0';
                when 169 => sda_i <= '0';
                when 170 => sda_i <= '0';
                when 171 => sda_i <= '0';
                when 172 => sda_i <= '0';
                when 173 => sda_i <= '0';
                when 174 => sda_i <= '0';
                when 175 => sda_i <= '0';
                when 176 => sda_i <= '0';
                when 177 => sda_i <= '0';
                when 178 => sda_i <= '0';
                when 179 => sda_i <= '0';
                when 180 => sda_i <= '1';
                when 181 => sda_i <= '1';
                when 182 => sda_i <= '1';
                when 183 => sda_i <= '1';
                when 184 => sda_i <= '1';
                when 185 => sda_i <= '1';
                when 186 => sda_i <= '1';
                when 187 => sda_i <= '1';
                when 188 => sda_i <= '1';
                when 189 => sda_i <= '1';
                when 190 => sda_i <= '1';
                when 191 => sda_i <= '1';
                when 192 => sda_i <= '1';
                when 193 => sda_i <= '1';
                when 194 => sda_i <= '1';
                when 195 => sda_i <= '1';
                when 196 => sda_i <= '1';
                when 197 => sda_i <= '1';
                when 198 => sda_i <= '1';
                when 199 => sda_i <= '1';
                when 200 => sda_i <= '1';
                when 201 => sda_i <= '1';
                when 202 => sda_i <= '1';
                when 203 => sda_i <= '1';
                when 204 => sda_i <= '1';
                when 205 => sda_i <= '1';
                when 206 => sda_i <= '1';
                when 207 => sda_i <= '1';
                when 208 => sda_i <= '1';
                when 209 => sda_i <= '1';
                when 210 => sda_i <= '1';
                when 211 => sda_i <= '1';
                when 212 => sda_i <= '1';
                when 213 => sda_i <= '0';
                when 214 => sda_i <= '0';
                when 215 => sda_i <= '0';
                when 216 => sda_i <= '0';
                when 217 => sda_i <= '0';
                when 218 => sda_i <= '0';
                when 219 => sda_i <= '0';
                when 220 => sda_i <= '0';
                when 221 => sda_i <= '0';
                when 222 => sda_i <= '0';
                when 223 => sda_i <= '0';
                when 224 => sda_i <= '0';
                when 225 => sda_i <= '0';
                when 226 => sda_i <= '0';
                when 227 => sda_i <= '0';
                when 228 => sda_i <= '0';
                when 229 => sda_i <= '0';
                when 230 => sda_i <= '0';
                when 231 => sda_i <= '0';
                when 232 => sda_i <= '0';
                when 233 => sda_i <= '0';
                when 234 => sda_i <= '0';
                when 235 => sda_i <= '0';
                when 236 => sda_i <= '0';
                when 237 => sda_i <= '0';
                when 238 => sda_i <= '0';
                when 239 => sda_i <= '0';
                when 240 => sda_i <= '0';
                when 241 => sda_i <= '0';
                when 242 => sda_i <= '0';
                when 243 => sda_i <= '0';
                when 244 => sda_i <= '0';
                when 245 => sda_i <= '0';
                when 246 => sda_i <= '0';
                when 247 => sda_i <= '0';
                when 248 => sda_i <= '0';
                when 249 => sda_i <= '0';
                when 250 => sda_i <= '0';
                when 251 => sda_i <= '0';
                when 252 => sda_i <= '0';
                when 253 => sda_i <= '0';
                when 254 => sda_i <= '0';
                when 255 => sda_i <= '0';
                when 256 => sda_i <= '0';
                when 257 => sda_i <= '0';
                when 258 => sda_i <= '0';
                when 259 => sda_i <= '0';
                when 260 => sda_i <= '0';
                when 261 => sda_i <= '0';
                when 262 => sda_i <= '0';
                when 263 => sda_i <= '0';
                when 264 => sda_i <= '0';
                when 265 => sda_i <= '0';
                when 266 => sda_i <= '0';
                when 267 => sda_i <= '0';
                when 268 => sda_i <= '0';
                when 269 => sda_i <= '0';
                when 270 => sda_i <= '0';
                when 271 => sda_i <= '0';
                when 272 => sda_i <= '0';
                when 273 => sda_i <= '0';
                when 274 => sda_i <= '0';
                when 275 => sda_i <= '0';
                when 276 => sda_i <= '0';
                when 277 => sda_i <= '0';
                when 278 => sda_i <= '0';
                when 279 => sda_i <= '0';
                when 280 => sda_i <= '0';
                when 281 => sda_i <= '0';
                when 282 => sda_i <= '0';
                when 283 => sda_i <= '0';
                when 284 => sda_i <= '0';
                when 285 => sda_i <= '0';
                when 286 => sda_i <= '0';
                when 287 => sda_i <= '0';
                when 288 => sda_i <= '0';
                when 289 => sda_i <= '0';
                when 290 => sda_i <= '0';
                when 291 => sda_i <= '0';
                when 292 => sda_i <= '0';
                when 293 => sda_i <= '0';
                when 294 => sda_i <= '0';
                when 295 => sda_i <= '0';
                when 296 => sda_i <= '0';
                when 297 => sda_i <= '0';
                when 298 => sda_i <= '0';
                when 299 => sda_i <= '0';
                when 300 => sda_i <= '0';
                when 301 => sda_i <= '0';
                when 302 => sda_i <= '0';
                when 303 => sda_i <= '0';
                when 304 => sda_i <= '0';
                when 305 => sda_i <= '0';
                when 306 => sda_i <= '0';
                when 307 => sda_i <= '0';
                when 308 => sda_i <= '0';
                when 309 => sda_i <= '0';
                when 310 => sda_i <= '0';
                when 311 => sda_i <= '0';
                when 312 => sda_i <= '0';
                when 313 => sda_i <= '0';
                when 314 => sda_i <= '0';
                when 315 => sda_i <= '0';
                when 316 => sda_i <= '0';
                when 317 => sda_i <= '0';
                when 318 => sda_i <= '0';
                when 319 => sda_i <= '0';
                when 320 => sda_i <= '0';
                when 321 => sda_i <= '0';
                when 322 => sda_i <= '1';
                when 323 => sda_i <= '1';
                when 324 => sda_i <= '0';
                when 325 => sda_i <= '0';
                when 326 => sda_i <= '0';
                when 327 => sda_i <= '0';
                when 328 => sda_i <= '0';
                when 329 => sda_i <= '0';
                when 330 => sda_i <= '0';
                when 331 => sda_i <= '0';
                when 332 => sda_i <= '0';
                when 333 => sda_i <= '0';
                when 334 => sda_i <= '0';
                when 335 => sda_i <= '0';
                when 336 => sda_i <= '0';
                when 337 => sda_i <= '0';
                when 338 => sda_i <= '0';
                when 339 => sda_i <= '0';
                when 340 => sda_i <= '0';
                when 341 => sda_i <= '0';
                when 342 => sda_i <= '0';
                when 343 => sda_i <= '0';
                when 344 => sda_i <= '0';
                when 345 => sda_i <= '0';
                when 346 => sda_i <= '0';
                when 347 => sda_i <= '0';
                when 348 => sda_i <= '0';
                when 349 => sda_i <= '0';
                when 350 => sda_i <= '0';
                when 351 => sda_i <= '0';
                when 352 => sda_i <= '0';
                when 353 => sda_i <= '0';
                when 354 => sda_i <= '0';
                when 355 => sda_i <= '0';
                when 356 => sda_i <= '0';
                when 357 => sda_i <= '0';
                when 358 => sda_i <= '0';
                when 359 => sda_i <= '0';
                when 360 => sda_i <= '0';
                when 361 => sda_i <= '0';
                when 362 => sda_i <= '0';
                when 363 => sda_i <= '0';
                when 364 => sda_i <= '0';
                when 365 => sda_i <= '0';
                when 366 => sda_i <= '0';
                when 367 => sda_i <= '0';
                when 368 => sda_i <= '0';
                when 369 => sda_i <= '0';
                when 370 => sda_i <= '0';
                when 371 => sda_i <= '0';
                when 372 => sda_i <= '0';
                when 373 => sda_i <= '0';
                when 374 => sda_i <= '0';
                when 375 => sda_i <= '0';
                when 376 => sda_i <= '0';
                when 377 => sda_i <= '0';
                when 378 => sda_i <= '0';
                when 379 => sda_i <= '0';
                when 380 => sda_i <= '0';
                when 381 => sda_i <= '0';
                when 382 => sda_i <= '0';
                when 383 => sda_i <= '0';
                when 384 => sda_i <= '0';
                when 385 => sda_i <= '0';
                when 386 => sda_i <= '0';
                when 387 => sda_i <= '0';
                when 388 => sda_i <= '0';
                when 389 => sda_i <= '0';
                when 390 => sda_i <= '0';
                when 391 => sda_i <= '0';
                when 392 => sda_i <= '0';
                when 393 => sda_i <= '0';
                when 394 => sda_i <= '0';
                when 395 => sda_i <= '0';
                when 396 => sda_i <= '0';
                when 397 => sda_i <= '0';
                when 398 => sda_i <= '0';
                when 399 => sda_i <= '0';
                when 400 => sda_i <= '0';
                when 401 => sda_i <= '0';
                when 402 => sda_i <= '0';
                when 403 => sda_i <= '0';
                when 404 => sda_i <= '0';
                when 405 => sda_i <= '0';
                when 406 => sda_i <= '0';
                when 407 => sda_i <= '0';
                when 408 => sda_i <= '0';
                when 409 => sda_i <= '0';
                when 410 => sda_i <= '0';
                when 411 => sda_i <= '0';
                when 412 => sda_i <= '0';
                when 413 => sda_i <= '0';
                when 414 => sda_i <= '0';
                when 415 => sda_i <= '0';
                when 416 => sda_i <= '0';
                when 417 => sda_i <= '0';
                when 418 => sda_i <= '0';
                when 419 => sda_i <= '0';
                when 420 => sda_i <= '0';
                when 421 => sda_i <= '0';
                when 422 => sda_i <= '0';
                when 423 => sda_i <= '0';
                when 424 => sda_i <= '0';
                when 425 => sda_i <= '0';
                when 426 => sda_i <= '0';
                when 427 => sda_i <= '0';
                when 428 => sda_i <= '0';
                when 429 => sda_i <= '0';
                when 430 => sda_i <= '1';
                when 431 => sda_i <= '1';
                when 432 => sda_i <= '0';
                when 433 => sda_i <= '0';
                when 434 => sda_i <= '0';
                when 435 => sda_i <= '0';
                when 436 => sda_i <= '0';
                when 437 => sda_i <= '0';
                when 438 => sda_i <= '0';
                when 439 => sda_i <= '0';
                when 440 => sda_i <= '0';
                when 441 => sda_i <= '0';
                when 442 => sda_i <= '0';
                when 443 => sda_i <= '0';
                when 444 => sda_i <= '0';
                when 445 => sda_i <= '0';
                when 446 => sda_i <= '0';
                when 447 => sda_i <= '0';
                when 448 => sda_i <= '0';
                when 449 => sda_i <= '0';
                when 450 => sda_i <= '0';
                when 451 => sda_i <= '0';
                when 452 => sda_i <= '0';
                when 453 => sda_i <= '0';
                when 454 => sda_i <= '0';
                when 455 => sda_i <= '0';
                when 456 => sda_i <= '0';
                when 457 => sda_i <= '0';
                when 458 => sda_i <= '0';
                when 459 => sda_i <= '0';
                when 460 => sda_i <= '0';
                when 461 => sda_i <= '0';
                when 462 => sda_i <= '0';
                when 463 => sda_i <= '0';
                when 464 => sda_i <= '0';
                when 465 => sda_i <= '0';
                when 466 => sda_i <= '0';
                when 467 => sda_i <= '0';
                when 468 => sda_i <= '0';
                when 469 => sda_i <= '0';
                when 470 => sda_i <= '0';
                when 471 => sda_i <= '0';
                when 472 => sda_i <= '0';
                when 473 => sda_i <= '0';
                when 474 => sda_i <= '0';
                when 475 => sda_i <= '0';
                when 476 => sda_i <= '0';
                when 477 => sda_i <= '0';
                when 478 => sda_i <= '0';
                when 479 => sda_i <= '0';
                when 480 => sda_i <= '0';
                when 481 => sda_i <= '0';
                when 482 => sda_i <= '0';
                when 483 => sda_i <= '0';
                when 484 => sda_i <= '0';
                when 485 => sda_i <= '0';
                when 486 => sda_i <= '0';
                when 487 => sda_i <= '0';
                when 488 => sda_i <= '0';
                when 489 => sda_i <= '0';
                when 490 => sda_i <= '0';
                when 491 => sda_i <= '0';
                when 492 => sda_i <= '0';
                when 493 => sda_i <= '0';
                when 494 => sda_i <= '0';
                when 495 => sda_i <= '0';
                when 496 => sda_i <= '0';
                when 497 => sda_i <= '0';
                when 498 => sda_i <= '0';
                when 499 => sda_i <= '0';
                when 500 => sda_i <= '0';
                when 501 => sda_i <= '0';
                when 502 => sda_i <= '0';
                when 503 => sda_i <= '0';
                when 504 => sda_i <= '0';
                when 505 => sda_i <= '0';
                when 506 => sda_i <= '0';
                when 507 => sda_i <= '0';
                when 508 => sda_i <= '0';
                when 509 => sda_i <= '0';
                when 510 => sda_i <= '0';
                when 511 => sda_i <= '0';
                when 512 => sda_i <= '0';
                when 513 => sda_i <= '0';
                when 514 => sda_i <= '0';
                when 515 => sda_i <= '0';
                when 516 => sda_i <= '0';
                when 517 => sda_i <= '0';
                when 518 => sda_i <= '0';
                when 519 => sda_i <= '0';
                when 520 => sda_i <= '0';
                when 521 => sda_i <= '0';
                when 522 => sda_i <= '0';
                when 523 => sda_i <= '0';
                when 524 => sda_i <= '0';
                when 525 => sda_i <= '0';
                when 526 => sda_i <= '0';
                when 527 => sda_i <= '0';
                when 528 => sda_i <= '0';
                when 529 => sda_i <= '0';
                when 530 => sda_i <= '0';
                when 531 => sda_i <= '0';
                when 532 => sda_i <= '0';
                when 533 => sda_i <= '0';
                when 534 => sda_i <= '0';
                when 535 => sda_i <= '0';
                when 536 => sda_i <= '0';
                when 537 => sda_i <= '0';
                when 538 => sda_i <= '1';
                when 539 => sda_i <= '1';
                when 540 => sda_i <= '0';
                when 541 => sda_i <= '0';
                when 542 => sda_i <= '0';
                when 543 => sda_i <= '0';
                when 544 => sda_i <= '0';
                when 545 => sda_i <= '0';
                when 546 => sda_i <= '0';
                when 547 => sda_i <= '0';
                when 548 => sda_i <= '0';
                when 549 => sda_i <= '0';
                when 550 => sda_i <= '0';
                when 551 => sda_i <= '0';
                when 552 => sda_i <= '0';
                when 553 => sda_i <= '0';
                when 554 => sda_i <= '0';
                when 555 => sda_i <= '0';
                when 556 => sda_i <= '0';
                when 557 => sda_i <= '0';
                when 558 => sda_i <= '0';
                when 559 => sda_i <= '0';
                when 560 => sda_i <= '0';
                when 561 => sda_i <= '0';
                when 562 => sda_i <= '0';
                when 563 => sda_i <= '0';
                when 564 => sda_i <= '0';
                when 565 => sda_i <= '0';
                when 566 => sda_i <= '0';
                when 567 => sda_i <= '0';
                when 568 => sda_i <= '0';
                when 569 => sda_i <= '0';
                when 570 => sda_i <= '0';
                when 571 => sda_i <= '0';
                when 572 => sda_i <= '0';
                when 573 => sda_i <= '0';
                when 574 => sda_i <= '0';
                when 575 => sda_i <= '0';
                when 576 => sda_i <= '0';
                when 577 => sda_i <= '0';
                when 578 => sda_i <= '0';
                when 579 => sda_i <= '0';
                when 580 => sda_i <= '0';
                when 581 => sda_i <= '0';
                when 582 => sda_i <= '0';
                when 583 => sda_i <= '0';
                when 584 => sda_i <= '0';
                when 585 => sda_i <= '0';
                when 586 => sda_i <= '0';
                when 587 => sda_i <= '0';
                when 588 => sda_i <= '0';
                when 589 => sda_i <= '0';
                when 590 => sda_i <= '0';
                when 591 => sda_i <= '0';
                when 592 => sda_i <= '0';
                when 593 => sda_i <= '0';
                when 594 => sda_i <= '0';
                when 595 => sda_i <= '0';
                when 596 => sda_i <= '0';
                when 597 => sda_i <= '0';
                when 598 => sda_i <= '0';
                when 599 => sda_i <= '0';
                when 600 => sda_i <= '0';
                when 601 => sda_i <= '0';
                when 602 => sda_i <= '0';
                when 603 => sda_i <= '0';
                when 604 => sda_i <= '0';
                when 605 => sda_i <= '0';
                when 606 => sda_i <= '0';
                when 607 => sda_i <= '0';
                when 608 => sda_i <= '0';
                when 609 => sda_i <= '0';
                when 610 => sda_i <= '0';
                when 611 => sda_i <= '0';
                when 612 => sda_i <= '0';
                when 613 => sda_i <= '0';
                when 614 => sda_i <= '0';
                when 615 => sda_i <= '0';
                when 616 => sda_i <= '0';
                when 617 => sda_i <= '0';
                when 618 => sda_i <= '0';
                when 619 => sda_i <= '0';
                when 620 => sda_i <= '0';
                when 621 => sda_i <= '0';
                when 622 => sda_i <= '0';
                when 623 => sda_i <= '0';
                when 624 => sda_i <= '0';
                when 625 => sda_i <= '0';
                when 626 => sda_i <= '0';
                when 627 => sda_i <= '0';
                when 628 => sda_i <= '0';
                when 629 => sda_i <= '0';
                when 630 => sda_i <= '0';
                when 631 => sda_i <= '0';
                when 632 => sda_i <= '0';
                when 633 => sda_i <= '0';
                when 634 => sda_i <= '0';
                when 635 => sda_i <= '0';
                when 636 => sda_i <= '0';
                when 637 => sda_i <= '0';
                when 638 => sda_i <= '0';
                when 639 => sda_i <= '0';
                when 640 => sda_i <= '0';
                when 641 => sda_i <= '0';
                when 642 => sda_i <= '0';
                when 643 => sda_i <= '0';
                when 644 => sda_i <= '0';
                when 645 => sda_i <= '0';
                when 646 => sda_i <= '1';
                when 647 => sda_i <= '1';
                when 648 => sda_i <= '0';
                when 649 => sda_i <= '0';
                when 650 => sda_i <= '0';
                when 651 => sda_i <= '0';
                when 652 => sda_i <= '0';
                when 653 => sda_i <= '0';
                when 654 => sda_i <= '0';
                when 655 => sda_i <= '0';
                when 656 => sda_i <= '0';
                when 657 => sda_i <= '0';
                when 658 => sda_i <= '0';
                when 659 => sda_i <= '0';
                when 660 => sda_i <= '0';
                when 661 => sda_i <= '0';
                when 662 => sda_i <= '0';
                when 663 => sda_i <= '0';
                when 664 => sda_i <= '0';
                when 665 => sda_i <= '0';
                when 666 => sda_i <= '0';
                when 667 => sda_i <= '0';
                when 668 => sda_i <= '0';
                when 669 => sda_i <= '0';
                when 670 => sda_i <= '0';
                when 671 => sda_i <= '0';
                when 672 => sda_i <= '0';
                when 673 => sda_i <= '0';
                when 674 => sda_i <= '0';
                when 675 => sda_i <= '0';
                when 676 => sda_i <= '0';
                when 677 => sda_i <= '0';
                when 678 => sda_i <= '0';
                when 679 => sda_i <= '0';
                when 680 => sda_i <= '0';
                when 681 => sda_i <= '0';
                when 682 => sda_i <= '0';
                when 683 => sda_i <= '0';
                when 684 => sda_i <= '0';
                when 685 => sda_i <= '0';
                when 686 => sda_i <= '0';
                when 687 => sda_i <= '0';
                when 688 => sda_i <= '0';
                when 689 => sda_i <= '0';
                when 690 => sda_i <= '0';
                when 691 => sda_i <= '0';
                when 692 => sda_i <= '0';
                when 693 => sda_i <= '0';
                when 694 => sda_i <= '0';
                when 695 => sda_i <= '0';
                when 696 => sda_i <= '0';
                when 697 => sda_i <= '0';
                when 698 => sda_i <= '0';
                when 699 => sda_i <= '0';
                when 700 => sda_i <= '0';
                when 701 => sda_i <= '0';
                when 702 => sda_i <= '0';
                when 703 => sda_i <= '0';
                when 704 => sda_i <= '0';
                when 705 => sda_i <= '0';
                when 706 => sda_i <= '1';
                when 707 => sda_i <= '1';
                when 708 => sda_i <= '1';
                when 709 => sda_i <= '1';
                when 710 => sda_i <= '1';
                when 711 => sda_i <= '1';
                when 712 => sda_i <= '1';
                when 713 => sda_i <= '1';
                when 714 => sda_i <= '1';
                when 715 => sda_i <= '1';
                when 716 => sda_i <= '1';
                when 717 => sda_i <= '0';
                when 718 => sda_i <= '0';
                when 719 => sda_i <= '0';
                when 720 => sda_i <= '0';
                when 721 => sda_i <= '0';
                when 722 => sda_i <= '0';
                when 723 => sda_i <= '0';
                when 724 => sda_i <= '0';
                when 725 => sda_i <= '0';
                when 726 => sda_i <= '0';
                when 727 => sda_i <= '0';
                when 728 => sda_i <= '0';
                when 729 => sda_i <= '0';
                when 730 => sda_i <= '1';
                when 731 => sda_i <= '1';
                when 732 => sda_i <= '1';
                when 733 => sda_i <= '1';
                when 734 => sda_i <= '1';
                when 735 => sda_i <= '1';
                when 736 => sda_i <= '1';
                when 737 => sda_i <= '1';
                when 738 => sda_i <= '1';
                when 739 => sda_i <= '1';
                when 740 => sda_i <= '1';
                when 741 => sda_i <= '0';
                when 742 => sda_i <= '0';
                when 743 => sda_i <= '0';
                when 744 => sda_i <= '0';
                when 745 => sda_i <= '0';
                when 746 => sda_i <= '0';
                when 747 => sda_i <= '0';
                when 748 => sda_i <= '0';
                when 749 => sda_i <= '0';
                when 750 => sda_i <= '0';
                when 751 => sda_i <= '0';
                when 752 => sda_i <= '0';
                when 753 => sda_i <= '0';
                when 754 => sda_i <= '1';
                when 755 => sda_i <= '1';
                when 756 => sda_i <= '0';
                when 757 => sda_i <= '0';
                when 758 => sda_i <= '0';
                when 759 => sda_i <= '0';
                when 760 => sda_i <= '0';
                when 761 => sda_i <= '0';
                when 762 => sda_i <= '0';
                when 763 => sda_i <= '0';
                when 764 => sda_i <= '0';
                when 765 => sda_i <= '0';
                when 766 => sda_i <= '0';
                when 767 => sda_i <= '0';
                when 768 => sda_i <= '0';
                when 769 => sda_i <= '0';
                when 770 => sda_i <= '0';
                when 771 => sda_i <= '0';
                when 772 => sda_i <= '0';
                when 773 => sda_i <= '0';
                when 774 => sda_i <= '0';
                when 775 => sda_i <= '0';
                when 776 => sda_i <= '0';
                when 777 => sda_i <= '0';
                when 778 => sda_i <= '0';
                when 779 => sda_i <= '0';
                when 780 => sda_i <= '0';
                when 781 => sda_i <= '0';
                when 782 => sda_i <= '0';
                when 783 => sda_i <= '0';
                when 784 => sda_i <= '0';
                when 785 => sda_i <= '0';
                when 786 => sda_i <= '0';
                when 787 => sda_i <= '0';
                when 788 => sda_i <= '0';
                when 789 => sda_i <= '0';
                when 790 => sda_i <= '0';
                when 791 => sda_i <= '0';
                when 792 => sda_i <= '0';
                when 793 => sda_i <= '0';
                when 794 => sda_i <= '0';
                when 795 => sda_i <= '0';
                when 796 => sda_i <= '0';
                when 797 => sda_i <= '0';
                when 798 => sda_i <= '0';
                when 799 => sda_i <= '0';
                when 800 => sda_i <= '0';
                when 801 => sda_i <= '0';
                when 802 => sda_i <= '0';
                when 803 => sda_i <= '0';
                when 804 => sda_i <= '0';
                when 805 => sda_i <= '0';
                when 806 => sda_i <= '0';
                when 807 => sda_i <= '0';
                when 808 => sda_i <= '0';
                when 809 => sda_i <= '0';
                when 810 => sda_i <= '0';
                when 811 => sda_i <= '0';
                when 812 => sda_i <= '0';
                when 813 => sda_i <= '0';
                when 814 => sda_i <= '0';
                when 815 => sda_i <= '0';
                when 816 => sda_i <= '0';
                when 817 => sda_i <= '0';
                when 818 => sda_i <= '0';
                when 819 => sda_i <= '0';
                when 820 => sda_i <= '0';
                when 821 => sda_i <= '0';
                when 822 => sda_i <= '0';
                when 823 => sda_i <= '0';
                when 824 => sda_i <= '0';
                when 825 => sda_i <= '0';
                when 826 => sda_i <= '0';
                when 827 => sda_i <= '0';
                when 828 => sda_i <= '0';
                when 829 => sda_i <= '0';
                when 830 => sda_i <= '0';
                when 831 => sda_i <= '0';
                when 832 => sda_i <= '0';
                when 833 => sda_i <= '0';
                when 834 => sda_i <= '0';
                when 835 => sda_i <= '0';
                when 836 => sda_i <= '0';
                when 837 => sda_i <= '0';
                when 838 => sda_i <= '0';
                when 839 => sda_i <= '0';
                when 840 => sda_i <= '0';
                when 841 => sda_i <= '0';
                when 842 => sda_i <= '0';
                when 843 => sda_i <= '0';
                when 844 => sda_i <= '0';
                when 845 => sda_i <= '0';
                when 846 => sda_i <= '0';
                when 847 => sda_i <= '0';
                when 848 => sda_i <= '0';
                when 849 => sda_i <= '0';
                when 850 => sda_i <= '0';
                when 851 => sda_i <= '0';
                when 852 => sda_i <= '0';
                when 853 => sda_i <= '0';
                when 854 => sda_i <= '0';
                when 855 => sda_i <= '0';
                when 856 => sda_i <= '0';
                when 857 => sda_i <= '0';
                when 858 => sda_i <= '0';
                when 859 => sda_i <= '0';
                when 860 => sda_i <= '0';
                when 861 => sda_i <= '0';
                when 862 => sda_i <= '1';
                when 863 => sda_i <= '1';
                when 864 => sda_i <= '0';
                when 865 => sda_i <= '0';
                when 866 => sda_i <= '0';
                when 867 => sda_i <= '0';
                when 868 => sda_i <= '0';
                when 869 => sda_i <= '0';
                when 870 => sda_i <= '0';
                when 871 => sda_i <= '0';
                when 872 => sda_i <= '0';
                when 873 => sda_i <= '0';
                when 874 => sda_i <= '0';
                when 875 => sda_i <= '0';
                when 876 => sda_i <= '0';
                when 877 => sda_i <= '0';
                when 878 => sda_i <= '0';
                when 879 => sda_i <= '0';
                when 880 => sda_i <= '0';
                when 881 => sda_i <= '0';
                when 882 => sda_i <= '0';
                when 883 => sda_i <= '0';
                when 884 => sda_i <= '0';
                when 885 => sda_i <= '0';
                when 886 => sda_i <= '0';
                when 887 => sda_i <= '0';
                when 888 => sda_i <= '0';
                when 889 => sda_i <= '0';
                when 890 => sda_i <= '0';
                when 891 => sda_i <= '0';
                when 892 => sda_i <= '0';
                when 893 => sda_i <= '0';
                when 894 => sda_i <= '0';
                when 895 => sda_i <= '0';
                when 896 => sda_i <= '0';
                when 897 => sda_i <= '0';
                when 898 => sda_i <= '0';
                when 899 => sda_i <= '0';
                when 900 => sda_i <= '0';
                when 901 => sda_i <= '0';
                when 902 => sda_i <= '0';
                when 903 => sda_i <= '0';
                when 904 => sda_i <= '0';
                when 905 => sda_i <= '0';
                when 906 => sda_i <= '0';
                when 907 => sda_i <= '0';
                when 908 => sda_i <= '0';
                when 909 => sda_i <= '0';
                when 910 => sda_i <= '0';
                when 911 => sda_i <= '0';
                when 912 => sda_i <= '0';
                when 913 => sda_i <= '0';
                when 914 => sda_i <= '0';
                when 915 => sda_i <= '0';
                when 916 => sda_i <= '0';
                when 917 => sda_i <= '0';
                when 918 => sda_i <= '0';
                when 919 => sda_i <= '0';
                when 920 => sda_i <= '0';
                when 921 => sda_i <= '0';
                when 922 => sda_i <= '0';
                when 923 => sda_i <= '0';
                when 924 => sda_i <= '0';
                when 925 => sda_i <= '0';
                when 926 => sda_i <= '0';
                when 927 => sda_i <= '0';
                when 928 => sda_i <= '0';
                when 929 => sda_i <= '0';
                when 930 => sda_i <= '0';
                when 931 => sda_i <= '0';
                when 932 => sda_i <= '0';
                when 933 => sda_i <= '0';
                when 934 => sda_i <= '0';
                when 935 => sda_i <= '0';
                when 936 => sda_i <= '0';
                when 937 => sda_i <= '0';
                when 938 => sda_i <= '0';
                when 939 => sda_i <= '0';
                when 940 => sda_i <= '0';
                when 941 => sda_i <= '0';
                when 942 => sda_i <= '0';
                when 943 => sda_i <= '0';
                when 944 => sda_i <= '0';
                when 945 => sda_i <= '0';
                when 946 => sda_i <= '0';
                when 947 => sda_i <= '0';
                when 948 => sda_i <= '0';
                when 949 => sda_i <= '0';
                when 950 => sda_i <= '0';
                when 951 => sda_i <= '0';
                when 952 => sda_i <= '0';
                when 953 => sda_i <= '0';
                when 954 => sda_i <= '0';
                when 955 => sda_i <= '0';
                when 956 => sda_i <= '0';
                when 957 => sda_i <= '0';
                when 958 => sda_i <= '0';
                when 959 => sda_i <= '0';
                when 960 => sda_i <= '0';
                when 961 => sda_i <= '0';
                when 962 => sda_i <= '0';
                when 963 => sda_i <= '0';
                when 964 => sda_i <= '0';
                when 965 => sda_i <= '0';
                when 966 => sda_i <= '0';
                when 967 => sda_i <= '0';
                when 968 => sda_i <= '0';
                when 969 => sda_i <= '0';
                when 970 => sda_i <= '1';
                when 971 => sda_i <= '1';
                when 972 => sda_i <= '0';
                when 973 => sda_i <= '0';
                when 974 => sda_i <= '0';
                when 975 => sda_i <= '0';
                when 976 => sda_i <= '0';
                when 977 => sda_i <= '0';
                when 978 => sda_i <= '0';
                when 979 => sda_i <= '0';
                when 980 => sda_i <= '0';
                when 981 => sda_i <= '0';
                when 982 => sda_i <= '0';
                when 983 => sda_i <= '0';
                when 984 => sda_i <= '0';
                when 985 => sda_i <= '0';
                when 986 => sda_i <= '0';
                when 987 => sda_i <= '0';
                when 988 => sda_i <= '0';
                when 989 => sda_i <= '0';
                when 990 => sda_i <= '0';
                when 991 => sda_i <= '0';
                when 992 => sda_i <= '0';
                when 993 => sda_i <= '0';
                when 994 => sda_i <= '0';
                when 995 => sda_i <= '0';
                when 996 => sda_i <= '0';
                when 997 => sda_i <= '0';
                when 998 => sda_i <= '0';
                when 999 => sda_i <= '0';
                when 1000 => sda_i <= '0';
                when 1001 => sda_i <= '0';
                when 1002 => sda_i <= '0';
                when 1003 => sda_i <= '0';
                when 1004 => sda_i <= '0';
                when 1005 => sda_i <= '0';
                when 1006 => sda_i <= '0';
                when 1007 => sda_i <= '0';
                when 1008 => sda_i <= '0';
                when 1009 => sda_i <= '0';
                when 1010 => sda_i <= '0';
                when 1011 => sda_i <= '0';
                when 1012 => sda_i <= '0';
                when 1013 => sda_i <= '0';
                when 1014 => sda_i <= '0';
                when 1015 => sda_i <= '0';
                when 1016 => sda_i <= '0';
                when 1017 => sda_i <= '0';
                when 1018 => sda_i <= '0';
                when 1019 => sda_i <= '0';
                when 1020 => sda_i <= '0';
                when 1021 => sda_i <= '0';
                when 1022 => sda_i <= '0';
                when 1023 => sda_i <= '0';
                when 1024 => sda_i <= '0';
                when 1025 => sda_i <= '0';
                when 1026 => sda_i <= '0';
                when 1027 => sda_i <= '0';
                when 1028 => sda_i <= '0';
                when 1029 => sda_i <= '0';
                when 1030 => sda_i <= '0';
                when 1031 => sda_i <= '0';
                when 1032 => sda_i <= '0';
                when 1033 => sda_i <= '0';
                when 1034 => sda_i <= '0';
                when 1035 => sda_i <= '0';
                when 1036 => sda_i <= '0';
                when 1037 => sda_i <= '0';
                when 1038 => sda_i <= '0';
                when 1039 => sda_i <= '0';
                when 1040 => sda_i <= '0';
                when 1041 => sda_i <= '0';
                when 1042 => sda_i <= '0';
                when 1043 => sda_i <= '0';
                when 1044 => sda_i <= '0';
                when 1045 => sda_i <= '0';
                when 1046 => sda_i <= '0';
                when 1047 => sda_i <= '0';
                when 1048 => sda_i <= '0';
                when 1049 => sda_i <= '0';
                when 1050 => sda_i <= '0';
                when 1051 => sda_i <= '0';
                when 1052 => sda_i <= '0';
                when 1053 => sda_i <= '0';
                when 1054 => sda_i <= '0';
                when 1055 => sda_i <= '0';
                when 1056 => sda_i <= '0';
                when 1057 => sda_i <= '0';
                when 1058 => sda_i <= '0';
                when 1059 => sda_i <= '0';
                when 1060 => sda_i <= '0';
                when 1061 => sda_i <= '0';
                when 1062 => sda_i <= '0';
                when 1063 => sda_i <= '0';
                when 1064 => sda_i <= '0';
                when 1065 => sda_i <= '0';
                when 1066 => sda_i <= '0';
                when 1067 => sda_i <= '0';
                when 1068 => sda_i <= '0';
                when 1069 => sda_i <= '0';
                when 1070 => sda_i <= '0';
                when 1071 => sda_i <= '0';
                when 1072 => sda_i <= '0';
                when 1073 => sda_i <= '0';
                when 1074 => sda_i <= '0';
                when 1075 => sda_i <= '0';
                when 1076 => sda_i <= '0';
                when 1077 => sda_i <= '0';
                when 1078 => sda_i <= '1';
                when 1079 => sda_i <= '1';
                when 1080 => sda_i <= '0';
                when 1081 => sda_i <= '0';
                when 1082 => sda_i <= '0';
                when 1083 => sda_i <= '0';
                when 1084 => sda_i <= '0';
                when 1085 => sda_i <= '0';
                when 1086 => sda_i <= '0';
                when 1087 => sda_i <= '0';
                when 1088 => sda_i <= '0';
                when 1089 => sda_i <= '0';
                when 1090 => sda_i <= '0';
                when 1091 => sda_i <= '0';
                when 1092 => sda_i <= '0';
                when 1093 => sda_i <= '0';
                when 1094 => sda_i <= '0';
                when 1095 => sda_i <= '0';
                when 1096 => sda_i <= '0';
                when 1097 => sda_i <= '0';
                when 1098 => sda_i <= '0';
                when 1099 => sda_i <= '0';
                when 1100 => sda_i <= '0';
                when 1101 => sda_i <= '0';
                when 1102 => sda_i <= '0';
                when 1103 => sda_i <= '0';
                when 1104 => sda_i <= '0';
                when 1105 => sda_i <= '0';
                when 1106 => sda_i <= '0';
                when 1107 => sda_i <= '0';
                when 1108 => sda_i <= '0';
                when 1109 => sda_i <= '0';
                when 1110 => sda_i <= '0';
                when 1111 => sda_i <= '0';
                when 1112 => sda_i <= '0';
                when 1113 => sda_i <= '0';
                when 1114 => sda_i <= '0';
                when 1115 => sda_i <= '0';
                when 1116 => sda_i <= '0';
                when 1117 => sda_i <= '0';
                when 1118 => sda_i <= '0';
                when 1119 => sda_i <= '0';
                when 1120 => sda_i <= '0';
                when 1121 => sda_i <= '0';
                when 1122 => sda_i <= '0';
                when 1123 => sda_i <= '0';
                when 1124 => sda_i <= '0';
                when 1125 => sda_i <= '0';
                when 1126 => sda_i <= '0';
                when 1127 => sda_i <= '0';
                when 1128 => sda_i <= '0';
                when 1129 => sda_i <= '0';
                when 1130 => sda_i <= '0';
                when 1131 => sda_i <= '0';
                when 1132 => sda_i <= '0';
                when 1133 => sda_i <= '0';
                when 1134 => sda_i <= '0';
                when 1135 => sda_i <= '0';
                when 1136 => sda_i <= '0';
                when 1137 => sda_i <= '0';
                when 1138 => sda_i <= '0';
                when 1139 => sda_i <= '0';
                when 1140 => sda_i <= '0';
                when 1141 => sda_i <= '0';
                when 1142 => sda_i <= '0';
                when 1143 => sda_i <= '0';
                when 1144 => sda_i <= '0';
                when 1145 => sda_i <= '0';
                when 1146 => sda_i <= '0';
                when 1147 => sda_i <= '0';
                when 1148 => sda_i <= '0';
                when 1149 => sda_i <= '0';
                when 1150 => sda_i <= '0';
                when 1151 => sda_i <= '0';
                when 1152 => sda_i <= '0';
                when 1153 => sda_i <= '0';
                when 1154 => sda_i <= '0';
                when 1155 => sda_i <= '0';
                when 1156 => sda_i <= '0';
                when 1157 => sda_i <= '0';
                when 1158 => sda_i <= '0';
                when 1159 => sda_i <= '0';
                when 1160 => sda_i <= '0';
                when 1161 => sda_i <= '0';
                when 1162 => sda_i <= '1';
                when 1163 => sda_i <= '1';
                when 1164 => sda_i <= '1';
                when 1165 => sda_i <= '1';
                when 1166 => sda_i <= '1';
                when 1167 => sda_i <= '1';
                when 1168 => sda_i <= '1';
                when 1169 => sda_i <= '1';
                when 1170 => sda_i <= '1';
                when 1171 => sda_i <= '1';
                when 1172 => sda_i <= '1';
                when 1173 => sda_i <= '0';
                when 1174 => sda_i <= '0';
                when 1175 => sda_i <= '0';
                when 1176 => sda_i <= '0';
                when 1177 => sda_i <= '0';
                when 1178 => sda_i <= '0';
                when 1179 => sda_i <= '0';
                when 1180 => sda_i <= '0';
                when 1181 => sda_i <= '0';
                when 1182 => sda_i <= '0';
                when 1183 => sda_i <= '0';
                when 1184 => sda_i <= '0';
                when 1185 => sda_i <= '0';
                when 1186 => sda_i <= '1';
                when 1187 => sda_i <= '1';
                when 1188 => sda_i <= '0';
                when 1189 => sda_i <= '0';
                when 1190 => sda_i <= '0';
                when 1191 => sda_i <= '0';
                when 1192 => sda_i <= '0';
                when 1193 => sda_i <= '0';
                when 1194 => sda_i <= '0';
                when 1195 => sda_i <= '0';
                when 1196 => sda_i <= '0';
                when 1197 => sda_i <= '0';
                when 1198 => sda_i <= '0';
                when 1199 => sda_i <= '0';
                when 1200 => sda_i <= '0';
                when 1201 => sda_i <= '0';
                when 1202 => sda_i <= '0';
                when 1203 => sda_i <= '0';
                when 1204 => sda_i <= '0';
                when 1205 => sda_i <= '0';
                when 1206 => sda_i <= '0';
                when 1207 => sda_i <= '0';
                when 1208 => sda_i <= '0';
                when 1209 => sda_i <= '0';
                when 1210 => sda_i <= '0';
                when 1211 => sda_i <= '0';
                when 1212 => sda_i <= '0';
                when 1213 => sda_i <= '0';
                when 1214 => sda_i <= '0';
                when 1215 => sda_i <= '0';
                when 1216 => sda_i <= '0';
                when 1217 => sda_i <= '0';
                when 1218 => sda_i <= '0';
                when 1219 => sda_i <= '0';
                when 1220 => sda_i <= '0';
                when 1221 => sda_i <= '0';
                when 1222 => sda_i <= '0';
                when 1223 => sda_i <= '0';
                when 1224 => sda_i <= '0';
                when 1225 => sda_i <= '0';
                when 1226 => sda_i <= '0';
                when 1227 => sda_i <= '0';
                when 1228 => sda_i <= '0';
                when 1229 => sda_i <= '0';
                when 1230 => sda_i <= '0';
                when 1231 => sda_i <= '0';
                when 1232 => sda_i <= '0';
                when 1233 => sda_i <= '0';
                when 1234 => sda_i <= '0';
                when 1235 => sda_i <= '0';
                when 1236 => sda_i <= '0';
                when 1237 => sda_i <= '0';
                when 1238 => sda_i <= '0';
                when 1239 => sda_i <= '0';
                when 1240 => sda_i <= '0';
                when 1241 => sda_i <= '0';
                when 1242 => sda_i <= '0';
                when 1243 => sda_i <= '0';
                when 1244 => sda_i <= '0';
                when 1245 => sda_i <= '0';
                when 1246 => sda_i <= '0';
                when 1247 => sda_i <= '0';
                when 1248 => sda_i <= '0';
                when 1249 => sda_i <= '0';
                when 1250 => sda_i <= '0';
                when 1251 => sda_i <= '0';
                when 1252 => sda_i <= '0';
                when 1253 => sda_i <= '0';
                when 1254 => sda_i <= '0';
                when 1255 => sda_i <= '0';
                when 1256 => sda_i <= '0';
                when 1257 => sda_i <= '0';
                when 1258 => sda_i <= '0';
                when 1259 => sda_i <= '0';
                when 1260 => sda_i <= '0';
                when 1261 => sda_i <= '0';
                when 1262 => sda_i <= '0';
                when 1263 => sda_i <= '0';
                when 1264 => sda_i <= '0';
                when 1265 => sda_i <= '0';
                when 1266 => sda_i <= '0';
                when 1267 => sda_i <= '0';
                when 1268 => sda_i <= '0';
                when 1269 => sda_i <= '0';
                when 1270 => sda_i <= '0';
                when 1271 => sda_i <= '0';
                when 1272 => sda_i <= '0';
                when 1273 => sda_i <= '0';
                when 1274 => sda_i <= '0';
                when 1275 => sda_i <= '0';
                when 1276 => sda_i <= '0';
                when 1277 => sda_i <= '0';
                when 1278 => sda_i <= '0';
                when 1279 => sda_i <= '0';
                when 1280 => sda_i <= '0';
                when 1281 => sda_i <= '0';
                when 1282 => sda_i <= '0';
                when 1283 => sda_i <= '0';
                when 1284 => sda_i <= '0';
                when 1285 => sda_i <= '0';
                when 1286 => sda_i <= '0';
                when 1287 => sda_i <= '0';
                when 1288 => sda_i <= '0';
                when 1289 => sda_i <= '0';
                when 1290 => sda_i <= '0';
                when 1291 => sda_i <= '0';
                when 1292 => sda_i <= '0';
                when 1293 => sda_i <= '0';
                when 1294 => sda_i <= '1';
                when 1295 => sda_i <= '1';
                when 1296 => sda_i <= '0';
                when 1297 => sda_i <= '0';
                when 1298 => sda_i <= '0';
                when 1299 => sda_i <= '0';
                when 1300 => sda_i <= '0';
                when 1301 => sda_i <= '0';
                when 1302 => sda_i <= '0';
                when 1303 => sda_i <= '0';
                when 1304 => sda_i <= '0';
                when 1305 => sda_i <= '0';
                when 1306 => sda_i <= '0';
                when 1307 => sda_i <= '0';
                when 1308 => sda_i <= '0';
                when 1309 => sda_i <= '0';
                when 1310 => sda_i <= '0';
                when 1311 => sda_i <= '0';
                when 1312 => sda_i <= '0';
                when 1313 => sda_i <= '0';
                when 1314 => sda_i <= '0';
                when 1315 => sda_i <= '0';
                when 1316 => sda_i <= '0';
                when 1317 => sda_i <= '0';
                when 1318 => sda_i <= '0';
                when 1319 => sda_i <= '0';
                when 1320 => sda_i <= '0';
                when 1321 => sda_i <= '0';
                when 1322 => sda_i <= '0';
                when 1323 => sda_i <= '0';
                when 1324 => sda_i <= '0';
                when 1325 => sda_i <= '0';
                when 1326 => sda_i <= '0';
                when 1327 => sda_i <= '0';
                when 1328 => sda_i <= '0';
                when 1329 => sda_i <= '0';
                when 1330 => sda_i <= '0';
                when 1331 => sda_i <= '0';
                when 1332 => sda_i <= '0';
                when 1333 => sda_i <= '0';
                when 1334 => sda_i <= '0';
                when 1335 => sda_i <= '0';
                when 1336 => sda_i <= '0';
                when 1337 => sda_i <= '0';
                when 1338 => sda_i <= '0';
                when 1339 => sda_i <= '0';
                when 1340 => sda_i <= '0';
                when 1341 => sda_i <= '0';
                when 1342 => sda_i <= '0';
                when 1343 => sda_i <= '0';
                when 1344 => sda_i <= '0';
                when 1345 => sda_i <= '0';
                when 1346 => sda_i <= '0';
                when 1347 => sda_i <= '0';
                when 1348 => sda_i <= '0';
                when 1349 => sda_i <= '0';
                when 1350 => sda_i <= '0';
                when 1351 => sda_i <= '0';
                when 1352 => sda_i <= '0';
                when 1353 => sda_i <= '0';
                when 1354 => sda_i <= '0';
                when 1355 => sda_i <= '0';
                when 1356 => sda_i <= '0';
                when 1357 => sda_i <= '0';
                when 1358 => sda_i <= '0';
                when 1359 => sda_i <= '0';
                when 1360 => sda_i <= '0';
                when 1361 => sda_i <= '0';
                when 1362 => sda_i <= '0';
                when 1363 => sda_i <= '0';
                when 1364 => sda_i <= '0';
                when 1365 => sda_i <= '0';
                when 1366 => sda_i <= '0';
                when 1367 => sda_i <= '0';
                when 1368 => sda_i <= '0';
                when 1369 => sda_i <= '0';
                when 1370 => sda_i <= '0';
                when 1371 => sda_i <= '0';
                when 1372 => sda_i <= '0';
                when 1373 => sda_i <= '0';
                when 1374 => sda_i <= '0';
                when 1375 => sda_i <= '0';
                when 1376 => sda_i <= '0';
                when 1377 => sda_i <= '0';
                when 1378 => sda_i <= '0';
                when 1379 => sda_i <= '0';
                when 1380 => sda_i <= '0';
                when 1381 => sda_i <= '0';
                when 1382 => sda_i <= '0';
                when 1383 => sda_i <= '0';
                when 1384 => sda_i <= '0';
                when 1385 => sda_i <= '0';
                when 1386 => sda_i <= '0';
                when 1387 => sda_i <= '0';
                when 1388 => sda_i <= '0';
                when 1389 => sda_i <= '0';
                when 1390 => sda_i <= '0';
                when 1391 => sda_i <= '0';
                when 1392 => sda_i <= '0';
                when 1393 => sda_i <= '0';
                when 1394 => sda_i <= '0';
                when 1395 => sda_i <= '0';
                when 1396 => sda_i <= '0';
                when 1397 => sda_i <= '0';
                when 1398 => sda_i <= '0';
                when 1399 => sda_i <= '0';
                when 1400 => sda_i <= '0';
                when 1401 => sda_i <= '0';
                when 1402 => sda_i <= '1';
                when 1403 => sda_i <= '1';
                when 1404 => sda_i <= '0';
                when 1405 => sda_i <= '0';
                when 1406 => sda_i <= '0';
                when 1407 => sda_i <= '0';
                when 1408 => sda_i <= '0';
                when 1409 => sda_i <= '0';
                when 1410 => sda_i <= '0';
                when 1411 => sda_i <= '0';
                when 1412 => sda_i <= '0';
                when 1413 => sda_i <= '0';
                when 1414 => sda_i <= '0';
                when 1415 => sda_i <= '0';
                when 1416 => sda_i <= '0';
                when 1417 => sda_i <= '0';
                when 1418 => sda_i <= '0';
                when 1419 => sda_i <= '0';
                when 1420 => sda_i <= '0';
                when 1421 => sda_i <= '0';
                when 1422 => sda_i <= '0';
                when 1423 => sda_i <= '0';
                when 1424 => sda_i <= '0';
                when 1425 => sda_i <= '0';
                when 1426 => sda_i <= '0';
                when 1427 => sda_i <= '0';
                when 1428 => sda_i <= '0';
                when 1429 => sda_i <= '0';
                when 1430 => sda_i <= '0';
                when 1431 => sda_i <= '0';
                when 1432 => sda_i <= '0';
                when 1433 => sda_i <= '0';
                when 1434 => sda_i <= '0';
                when 1435 => sda_i <= '0';
                when 1436 => sda_i <= '0';
                when 1437 => sda_i <= '0';
                when 1438 => sda_i <= '0';
                when 1439 => sda_i <= '0';
                when 1440 => sda_i <= '0';
                when 1441 => sda_i <= '0';
                when 1442 => sda_i <= '0';
                when 1443 => sda_i <= '0';
                when 1444 => sda_i <= '0';
                when 1445 => sda_i <= '0';
                when 1446 => sda_i <= '0';
                when 1447 => sda_i <= '0';
                when 1448 => sda_i <= '0';
                when 1449 => sda_i <= '0';
                when 1450 => sda_i <= '0';
                when 1451 => sda_i <= '0';
                when 1452 => sda_i <= '0';
                when 1453 => sda_i <= '0';
                when 1454 => sda_i <= '0';
                when 1455 => sda_i <= '0';
                when 1456 => sda_i <= '0';
                when 1457 => sda_i <= '0';
                when 1458 => sda_i <= '0';
                when 1459 => sda_i <= '0';
                when 1460 => sda_i <= '0';
                when 1461 => sda_i <= '0';
                when 1462 => sda_i <= '0';
                when 1463 => sda_i <= '0';
                when 1464 => sda_i <= '0';
                when 1465 => sda_i <= '0';
                when 1466 => sda_i <= '0';
                when 1467 => sda_i <= '0';
                when 1468 => sda_i <= '0';
                when 1469 => sda_i <= '0';
                when 1470 => sda_i <= '0';
                when 1471 => sda_i <= '0';
                when 1472 => sda_i <= '0';
                when 1473 => sda_i <= '0';
                when 1474 => sda_i <= '0';
                when 1475 => sda_i <= '0';
                when 1476 => sda_i <= '0';
                when 1477 => sda_i <= '0';
                when 1478 => sda_i <= '0';
                when 1479 => sda_i <= '0';
                when 1480 => sda_i <= '0';
                when 1481 => sda_i <= '0';
                when 1482 => sda_i <= '0';
                when 1483 => sda_i <= '0';
                when 1484 => sda_i <= '0';
                when 1485 => sda_i <= '0';
                when 1486 => sda_i <= '0';
                when 1487 => sda_i <= '0';
                when 1488 => sda_i <= '0';
                when 1489 => sda_i <= '0';
                when 1490 => sda_i <= '0';
                when 1491 => sda_i <= '0';
                when 1492 => sda_i <= '0';
                when 1493 => sda_i <= '0';
                when 1494 => sda_i <= '0';
                when 1495 => sda_i <= '0';
                when 1496 => sda_i <= '0';
                when 1497 => sda_i <= '0';
                when 1498 => sda_i <= '0';
                when 1499 => sda_i <= '0';
                when 1500 => sda_i <= '0';
                when 1501 => sda_i <= '0';
                when 1502 => sda_i <= '0';
                when 1503 => sda_i <= '0';
                when 1504 => sda_i <= '0';
                when 1505 => sda_i <= '0';
                when 1506 => sda_i <= '0';
                when 1507 => sda_i <= '0';
                when 1508 => sda_i <= '0';
                when 1509 => sda_i <= '0';
                when 1510 => sda_i <= '1';
                when 1511 => sda_i <= '1';
                when 1512 => sda_i <= '0';
                when 1513 => sda_i <= '0';
                when 1514 => sda_i <= '0';
                when 1515 => sda_i <= '0';
                when 1516 => sda_i <= '0';
                when 1517 => sda_i <= '0';
                when 1518 => sda_i <= '0';
                when 1519 => sda_i <= '0';
                when 1520 => sda_i <= '0';
                when 1521 => sda_i <= '0';
                when 1522 => sda_i <= '0';
                when 1523 => sda_i <= '0';
                when 1524 => sda_i <= '0';
                when 1525 => sda_i <= '0';
                when 1526 => sda_i <= '0';
                when 1527 => sda_i <= '0';
                when 1528 => sda_i <= '0';
                when 1529 => sda_i <= '0';
                when 1530 => sda_i <= '0';
                when 1531 => sda_i <= '0';
                when 1532 => sda_i <= '0';
                when 1533 => sda_i <= '0';
                when 1534 => sda_i <= '0';
                when 1535 => sda_i <= '0';
                when 1536 => sda_i <= '0';
                when 1537 => sda_i <= '0';
                when 1538 => sda_i <= '0';
                when 1539 => sda_i <= '0';
                when 1540 => sda_i <= '0';
                when 1541 => sda_i <= '0';
                when 1542 => sda_i <= '0';
                when 1543 => sda_i <= '0';
                when 1544 => sda_i <= '0';
                when 1545 => sda_i <= '0';
                when 1546 => sda_i <= '0';
                when 1547 => sda_i <= '0';
                when 1548 => sda_i <= '0';
                when 1549 => sda_i <= '0';
                when 1550 => sda_i <= '0';
                when 1551 => sda_i <= '0';
                when 1552 => sda_i <= '0';
                when 1553 => sda_i <= '0';
                when 1554 => sda_i <= '0';
                when 1555 => sda_i <= '0';
                when 1556 => sda_i <= '0';
                when 1557 => sda_i <= '0';
                when 1558 => sda_i <= '0';
                when 1559 => sda_i <= '0';
                when 1560 => sda_i <= '0';
                when 1561 => sda_i <= '0';
                when 1562 => sda_i <= '0';
                when 1563 => sda_i <= '0';
                when 1564 => sda_i <= '0';
                when 1565 => sda_i <= '0';
                when 1566 => sda_i <= '0';
                when 1567 => sda_i <= '0';
                when 1568 => sda_i <= '0';
                when 1569 => sda_i <= '0';
                when 1570 => sda_i <= '0';
                when 1571 => sda_i <= '0';
                when 1572 => sda_i <= '0';
                when 1573 => sda_i <= '0';
                when 1574 => sda_i <= '0';
                when 1575 => sda_i <= '0';
                when 1576 => sda_i <= '0';
                when 1577 => sda_i <= '0';
                when 1578 => sda_i <= '0';
                when 1579 => sda_i <= '0';
                when 1580 => sda_i <= '0';
                when 1581 => sda_i <= '0';
                when 1582 => sda_i <= '0';
                when 1583 => sda_i <= '0';
                when 1584 => sda_i <= '0';
                when 1585 => sda_i <= '0';
                when 1586 => sda_i <= '0';
                when 1587 => sda_i <= '0';
                when 1588 => sda_i <= '0';
                when 1589 => sda_i <= '0';
                when 1590 => sda_i <= '0';
                when 1591 => sda_i <= '0';
                when 1592 => sda_i <= '0';
                when 1593 => sda_i <= '0';
                when 1594 => sda_i <= '0';
                when 1595 => sda_i <= '0';
                when 1596 => sda_i <= '0';
                when 1597 => sda_i <= '0';
                when 1598 => sda_i <= '0';
                when 1599 => sda_i <= '0';
                when 1600 => sda_i <= '0';
                when 1601 => sda_i <= '0';
                when 1602 => sda_i <= '0';
                when 1603 => sda_i <= '0';
                when 1604 => sda_i <= '0';
                when 1605 => sda_i <= '0';
                when 1606 => sda_i <= '0';
                when 1607 => sda_i <= '0';
                when 1608 => sda_i <= '0';
                when 1609 => sda_i <= '0';
                when 1610 => sda_i <= '0';
                when 1611 => sda_i <= '0';
                when 1612 => sda_i <= '0';
                when 1613 => sda_i <= '0';
                when 1614 => sda_i <= '0';
                when 1615 => sda_i <= '0';
                when 1616 => sda_i <= '0';
                when 1617 => sda_i <= '0';
                when 1618 => sda_i <= '1';
                when 1619 => sda_i <= '1';
                when 1620 => sda_i <= '0';
                when 1621 => sda_i <= '0';
                when 1622 => sda_i <= '0';
                when 1623 => sda_i <= '0';
                when 1624 => sda_i <= '0';
                when 1625 => sda_i <= '0';
                when 1626 => sda_i <= '0';
                when 1627 => sda_i <= '0';
                when 1628 => sda_i <= '0';
                when 1629 => sda_i <= '0';
                when 1630 => sda_i <= '0';
                when 1631 => sda_i <= '0';
                when 1632 => sda_i <= '0';
                when 1633 => sda_i <= '0';
                when 1634 => sda_i <= '0';
                when 1635 => sda_i <= '0';
                when 1636 => sda_i <= '0';
                when 1637 => sda_i <= '0';
                when 1638 => sda_i <= '0';
                when 1639 => sda_i <= '0';
                when 1640 => sda_i <= '0';
                when 1641 => sda_i <= '0';
                when 1642 => sda_i <= '0';
                when 1643 => sda_i <= '0';
                when 1644 => sda_i <= '0';
                when 1645 => sda_i <= '0';
                when 1646 => sda_i <= '0';
                when 1647 => sda_i <= '0';
                when 1648 => sda_i <= '0';
                when 1649 => sda_i <= '0';
                when 1650 => sda_i <= '0';
                when 1651 => sda_i <= '0';
                when 1652 => sda_i <= '0';
                when 1653 => sda_i <= '0';
                when 1654 => sda_i <= '0';
                when 1655 => sda_i <= '0';
                when 1656 => sda_i <= '0';
                when 1657 => sda_i <= '0';
                when 1658 => sda_i <= '0';
                when 1659 => sda_i <= '0';
                when 1660 => sda_i <= '0';
                when 1661 => sda_i <= '0';
                when 1662 => sda_i <= '0';
                when 1663 => sda_i <= '0';
                when 1664 => sda_i <= '0';
                when 1665 => sda_i <= '0';
                when 1666 => sda_i <= '0';
                when 1667 => sda_i <= '0';
                when 1668 => sda_i <= '0';
                when 1669 => sda_i <= '0';
                when 1670 => sda_i <= '0';
                when 1671 => sda_i <= '0';
                when 1672 => sda_i <= '0';
                when 1673 => sda_i <= '0';
                when 1674 => sda_i <= '0';
                when 1675 => sda_i <= '0';
                when 1676 => sda_i <= '0';
                when 1677 => sda_i <= '0';
                when 1678 => sda_i <= '0';
                when 1679 => sda_i <= '0';
                when 1680 => sda_i <= '0';
                when 1681 => sda_i <= '0';
                when 1682 => sda_i <= '0';
                when 1683 => sda_i <= '0';
                when 1684 => sda_i <= '0';
                when 1685 => sda_i <= '0';
                when 1686 => sda_i <= '0';
                when 1687 => sda_i <= '0';
                when 1688 => sda_i <= '0';
                when 1689 => sda_i <= '0';
                when 1690 => sda_i <= '0';
                when 1691 => sda_i <= '0';
                when 1692 => sda_i <= '0';
                when 1693 => sda_i <= '0';
                when 1694 => sda_i <= '0';
                when 1695 => sda_i <= '0';
                when 1696 => sda_i <= '0';
                when 1697 => sda_i <= '0';
                when 1698 => sda_i <= '0';
                when 1699 => sda_i <= '0';
                when 1700 => sda_i <= '0';
                when 1701 => sda_i <= '0';
                when 1702 => sda_i <= '0';
                when 1703 => sda_i <= '0';
                when 1704 => sda_i <= '0';
                when 1705 => sda_i <= '0';
                when 1706 => sda_i <= '0';
                when 1707 => sda_i <= '0';
                when 1708 => sda_i <= '0';
                when 1709 => sda_i <= '0';
                when 1710 => sda_i <= '0';
                when 1711 => sda_i <= '0';
                when 1712 => sda_i <= '0';
                when 1713 => sda_i <= '0';
                when 1714 => sda_i <= '0';
                when 1715 => sda_i <= '0';
                when 1716 => sda_i <= '0';
                when 1717 => sda_i <= '0';
                when 1718 => sda_i <= '0';
                when 1719 => sda_i <= '0';
                when 1720 => sda_i <= '0';
                when 1721 => sda_i <= '0';
                when 1722 => sda_i <= '0';
                when 1723 => sda_i <= '0';
                when 1724 => sda_i <= '0';
                when 1725 => sda_i <= '0';
                when 1726 => sda_i <= '1';
                when 1727 => sda_i <= '1';
                when 1728 => sda_i <= '0';
                when 1729 => sda_i <= '0';
                when 1730 => sda_i <= '0';
                when 1731 => sda_i <= '0';
                when 1732 => sda_i <= '0';
                when 1733 => sda_i <= '0';
                when 1734 => sda_i <= '0';
                when 1735 => sda_i <= '0';
                when 1736 => sda_i <= '0';
                when 1737 => sda_i <= '0';
                when 1738 => sda_i <= '0';
                when 1739 => sda_i <= '0';
                when 1740 => sda_i <= '0';
                when 1741 => sda_i <= '0';
                when 1742 => sda_i <= '0';
                when 1743 => sda_i <= '0';
                when 1744 => sda_i <= '0';
                when 1745 => sda_i <= '0';
                when 1746 => sda_i <= '0';
                when 1747 => sda_i <= '0';
                when 1748 => sda_i <= '0';
                when 1749 => sda_i <= '0';
                when 1750 => sda_i <= '0';
                when 1751 => sda_i <= '0';
                when 1752 => sda_i <= '0';
                when 1753 => sda_i <= '0';
                when 1754 => sda_i <= '0';
                when 1755 => sda_i <= '0';
                when 1756 => sda_i <= '0';
                when 1757 => sda_i <= '0';
                when 1758 => sda_i <= '0';
                when 1759 => sda_i <= '0';
                when 1760 => sda_i <= '0';
                when 1761 => sda_i <= '0';
                when 1762 => sda_i <= '0';
                when 1763 => sda_i <= '0';
                when 1764 => sda_i <= '0';
                when 1765 => sda_i <= '0';
                when 1766 => sda_i <= '0';
                when 1767 => sda_i <= '0';
                when 1768 => sda_i <= '0';
                when 1769 => sda_i <= '0';
                when 1770 => sda_i <= '0';
                when 1771 => sda_i <= '0';
                when 1772 => sda_i <= '0';
                when 1773 => sda_i <= '0';
                when 1774 => sda_i <= '0';
                when 1775 => sda_i <= '0';
                when 1776 => sda_i <= '0';
                when 1777 => sda_i <= '0';
                when 1778 => sda_i <= '0';
                when 1779 => sda_i <= '0';
                when 1780 => sda_i <= '0';
                when 1781 => sda_i <= '0';
                when 1782 => sda_i <= '0';
                when 1783 => sda_i <= '0';
                when 1784 => sda_i <= '0';
                when 1785 => sda_i <= '0';
                when 1786 => sda_i <= '0';
                when 1787 => sda_i <= '0';
                when 1788 => sda_i <= '0';
                when 1789 => sda_i <= '0';
                when 1790 => sda_i <= '0';
                when 1791 => sda_i <= '0';
                when 1792 => sda_i <= '0';
                when 1793 => sda_i <= '0';
                when 1794 => sda_i <= '0';
                when 1795 => sda_i <= '0';
                when 1796 => sda_i <= '0';
                when 1797 => sda_i <= '0';
                when 1798 => sda_i <= '0';
                when 1799 => sda_i <= '0';
                when 1800 => sda_i <= '0';
                when 1801 => sda_i <= '0';
                when 1802 => sda_i <= '0';
                when 1803 => sda_i <= '0';
                when 1804 => sda_i <= '0';
                when 1805 => sda_i <= '0';
                when 1806 => sda_i <= '0';
                when 1807 => sda_i <= '0';
                when 1808 => sda_i <= '0';
                when 1809 => sda_i <= '0';
                when 1810 => sda_i <= '0';
                when 1811 => sda_i <= '0';
                when 1812 => sda_i <= '0';
                when 1813 => sda_i <= '0';
                when 1814 => sda_i <= '0';
                when 1815 => sda_i <= '0';
                when 1816 => sda_i <= '0';
                when 1817 => sda_i <= '0';
                when 1818 => sda_i <= '0';
                when 1819 => sda_i <= '0';
                when 1820 => sda_i <= '0';
                when 1821 => sda_i <= '0';
                when 1822 => sda_i <= '0';
                when 1823 => sda_i <= '0';
                when 1824 => sda_i <= '0';
                when 1825 => sda_i <= '0';
                when 1826 => sda_i <= '0';
                when 1827 => sda_i <= '0';
                when 1828 => sda_i <= '0';
                when 1829 => sda_i <= '0';
                when 1830 => sda_i <= '0';
                when 1831 => sda_i <= '0';
                when 1832 => sda_i <= '0';
                when 1833 => sda_i <= '0';
                when 1834 => sda_i <= '1';
                when 1835 => sda_i <= '1';
                when 1836 => sda_i <= '0';
                when 1837 => sda_i <= '0';
                when 1838 => sda_i <= '0';
                when 1839 => sda_i <= '0';
                when 1840 => sda_i <= '0';
                when 1841 => sda_i <= '0';
                when 1842 => sda_i <= '0';
                when 1843 => sda_i <= '0';
                when 1844 => sda_i <= '0';
                when 1845 => sda_i <= '0';
                when 1846 => sda_i <= '0';
                when 1847 => sda_i <= '0';
                when 1848 => sda_i <= '0';
                when 1849 => sda_i <= '0';
                when 1850 => sda_i <= '0';
                when 1851 => sda_i <= '0';
                when 1852 => sda_i <= '0';
                when 1853 => sda_i <= '0';
                when 1854 => sda_i <= '0';
                when 1855 => sda_i <= '0';
                when 1856 => sda_i <= '0';
                when 1857 => sda_i <= '0';
                when 1858 => sda_i <= '0';
                when 1859 => sda_i <= '0';
                when 1860 => sda_i <= '0';
                when 1861 => sda_i <= '0';
                when 1862 => sda_i <= '0';
                when 1863 => sda_i <= '0';
                when 1864 => sda_i <= '0';
                when 1865 => sda_i <= '0';
                when 1866 => sda_i <= '0';
                when 1867 => sda_i <= '0';
                when 1868 => sda_i <= '0';
                when 1869 => sda_i <= '0';
                when 1870 => sda_i <= '0';
                when 1871 => sda_i <= '0';
                when 1872 => sda_i <= '0';
                when 1873 => sda_i <= '0';
                when 1874 => sda_i <= '0';
                when 1875 => sda_i <= '0';
                when 1876 => sda_i <= '0';
                when 1877 => sda_i <= '0';
                when 1878 => sda_i <= '0';
                when 1879 => sda_i <= '0';
                when 1880 => sda_i <= '0';
                when 1881 => sda_i <= '0';
                when 1882 => sda_i <= '0';
                when 1883 => sda_i <= '0';
                when 1884 => sda_i <= '0';
                when 1885 => sda_i <= '0';
                when 1886 => sda_i <= '0';
                when 1887 => sda_i <= '0';
                when 1888 => sda_i <= '0';
                when 1889 => sda_i <= '0';
                when 1890 => sda_i <= '0';
                when 1891 => sda_i <= '0';
                when 1892 => sda_i <= '0';
                when 1893 => sda_i <= '0';
                when 1894 => sda_i <= '0';
                when 1895 => sda_i <= '0';
                when 1896 => sda_i <= '0';
                when 1897 => sda_i <= '0';
                when 1898 => sda_i <= '0';
                when 1899 => sda_i <= '0';
                when 1900 => sda_i <= '0';
                when 1901 => sda_i <= '0';
                when 1902 => sda_i <= '0';
                when 1903 => sda_i <= '0';
                when 1904 => sda_i <= '0';
                when 1905 => sda_i <= '0';
                when 1906 => sda_i <= '0';
                when 1907 => sda_i <= '0';
                when 1908 => sda_i <= '0';
                when 1909 => sda_i <= '0';
                when 1910 => sda_i <= '0';
                when 1911 => sda_i <= '0';
                when 1912 => sda_i <= '0';
                when 1913 => sda_i <= '0';
                when 1914 => sda_i <= '0';
                when 1915 => sda_i <= '0';
                when 1916 => sda_i <= '0';
                when 1917 => sda_i <= '0';
                when 1918 => sda_i <= '0';
                when 1919 => sda_i <= '0';
                when 1920 => sda_i <= '0';
                when 1921 => sda_i <= '0';
                when 1922 => sda_i <= '0';
                when 1923 => sda_i <= '0';
                when 1924 => sda_i <= '0';
                when 1925 => sda_i <= '0';
                when 1926 => sda_i <= '0';
                when 1927 => sda_i <= '0';
                when 1928 => sda_i <= '0';
                when 1929 => sda_i <= '0';
                when 1930 => sda_i <= '0';
                when 1931 => sda_i <= '0';
                when 1932 => sda_i <= '0';
                when 1933 => sda_i <= '0';
                when 1934 => sda_i <= '0';
                when 1935 => sda_i <= '0';
                when 1936 => sda_i <= '0';
                when 1937 => sda_i <= '0';
                when 1938 => sda_i <= '0';
                when 1939 => sda_i <= '0';
                when 1940 => sda_i <= '0';
                when 1941 => sda_i <= '0';
                when 1942 => sda_i <= '1';
                when 1943 => sda_i <= '1';
                when 1944 => sda_i <= '0';
                when 1945 => sda_i <= '0';
                when 1946 => sda_i <= '0';
                when 1947 => sda_i <= '0';
                when 1948 => sda_i <= '0';
                when 1949 => sda_i <= '0';
                when 1950 => sda_i <= '0';
                when 1951 => sda_i <= '0';
                when 1952 => sda_i <= '0';
                when 1953 => sda_i <= '0';
                when 1954 => sda_i <= '0';
                when 1955 => sda_i <= '0';
                when 1956 => sda_i <= '0';
                when 1957 => sda_i <= '0';
                when 1958 => sda_i <= '0';
                when 1959 => sda_i <= '0';
                when 1960 => sda_i <= '0';
                when 1961 => sda_i <= '0';
                when 1962 => sda_i <= '0';
                when 1963 => sda_i <= '0';
                when 1964 => sda_i <= '0';
                when 1965 => sda_i <= '0';
                when 1966 => sda_i <= '0';
                when 1967 => sda_i <= '0';
                when 1968 => sda_i <= '0';
                when 1969 => sda_i <= '0';
                when 1970 => sda_i <= '0';
                when 1971 => sda_i <= '0';
                when 1972 => sda_i <= '0';
                when 1973 => sda_i <= '0';
                when 1974 => sda_i <= '0';
                when 1975 => sda_i <= '0';
                when 1976 => sda_i <= '0';
                when 1977 => sda_i <= '0';
                when 1978 => sda_i <= '0';
                when 1979 => sda_i <= '0';
                when 1980 => sda_i <= '0';
                when 1981 => sda_i <= '0';
                when 1982 => sda_i <= '0';
                when 1983 => sda_i <= '0';
                when 1984 => sda_i <= '0';
                when 1985 => sda_i <= '0';
                when 1986 => sda_i <= '0';
                when 1987 => sda_i <= '0';
                when 1988 => sda_i <= '0';
                when 1989 => sda_i <= '0';
                when 1990 => sda_i <= '0';
                when 1991 => sda_i <= '0';
                when 1992 => sda_i <= '0';
                when 1993 => sda_i <= '0';
                when 1994 => sda_i <= '0';
                when 1995 => sda_i <= '0';
                when 1996 => sda_i <= '0';
                when 1997 => sda_i <= '0';
                when 1998 => sda_i <= '0';
                when 1999 => sda_i <= '0';

                when 2000 => sda_i <= '0';
                when 2001 => sda_i <= '0';
                when 2002 => sda_i <= '0';
                when 2003 => sda_i <= '0';
                when 2004 => sda_i <= '0';
                when 2005 => sda_i <= '0';
                when 2006 => sda_i <= '0';
                when 2007 => sda_i <= '0';
                when 2008 => sda_i <= '0';
                when 2009 => sda_i <= '0';
                when 2010 => sda_i <= '0';
                when 2011 => sda_i <= '0';
                when 2012 => sda_i <= '0';
                when 2013 => sda_i <= '0';
                when 2014 => sda_i <= '0';
                when 2015 => sda_i <= '0';
                when 2016 => sda_i <= '0';
                when 2017 => sda_i <= '0';
                when 2018 => sda_i <= '0';
                when 2019 => sda_i <= '0';
                when 2020 => sda_i <= '0';
                when 2021 => sda_i <= '0';
                when 2022 => sda_i <= '0';
                when 2023 => sda_i <= '0';
                when 2024 => sda_i <= '0';
                when 2025 => sda_i <= '0';
                when 2026 => sda_i <= '0';
                when 2027 => sda_i <= '0';
                when 2028 => sda_i <= '0';
                when 2029 => sda_i <= '0';
                when 2030 => sda_i <= '0';
                when 2031 => sda_i <= '0';
                when 2032 => sda_i <= '0';
                when 2033 => sda_i <= '0';
                when 2034 => sda_i <= '0';
                when 2035 => sda_i <= '0';
                when 2036 => sda_i <= '0';
                when 2037 => sda_i <= '0';
                when 2038 => sda_i <= '0';
                when 2039 => sda_i <= '0';
                when 2040 => sda_i <= '0';
                when 2041 => sda_i <= '0';
                when 2042 => sda_i <= '0';
                when 2043 => sda_i <= '0';
                when 2044 => sda_i <= '0';
                when 2045 => sda_i <= '0';
                when 2046 => sda_i <= '0';
                when 2047 => sda_i <= '0';
                when 2048 => sda_i <= '0';
                when 2049 => sda_i <= '0';
                when 2050 => sda_i <= '1';
                when 2051 => sda_i <= '1';
                when 2052 => sda_i <= '0';
                when 2053 => sda_i <= '0';
                when 2054 => sda_i <= '0';
                when 2055 => sda_i <= '0';
                when 2056 => sda_i <= '0';
                when 2057 => sda_i <= '0';
                when 2058 => sda_i <= '0';
                when 2059 => sda_i <= '0';
                when 2060 => sda_i <= '0';
                when 2061 => sda_i <= '0';
                when 2062 => sda_i <= '0';
                when 2063 => sda_i <= '0';
                when 2064 => sda_i <= '0';
                when 2065 => sda_i <= '0';
                when 2066 => sda_i <= '0';
                when 2067 => sda_i <= '0';
                when 2068 => sda_i <= '0';
                when 2069 => sda_i <= '0';
                when 2070 => sda_i <= '0';
                when 2071 => sda_i <= '0';
                when 2072 => sda_i <= '0';
                when 2073 => sda_i <= '0';
                when 2074 => sda_i <= '0';
                when 2075 => sda_i <= '0';
                when 2076 => sda_i <= '0';
                when 2077 => sda_i <= '0';
                when 2078 => sda_i <= '0';
                when 2079 => sda_i <= '0';
                when 2080 => sda_i <= '0';
                when 2081 => sda_i <= '0';
                when 2082 => sda_i <= '0';
                when 2083 => sda_i <= '0';
                when 2084 => sda_i <= '0';
                when 2085 => sda_i <= '0';
                when 2086 => sda_i <= '0';
                when 2087 => sda_i <= '0';
                when 2088 => sda_i <= '0';
                when 2089 => sda_i <= '0';
                when 2090 => sda_i <= '0';
                when 2091 => sda_i <= '0';
                when 2092 => sda_i <= '0';
                when 2093 => sda_i <= '0';
                when 2094 => sda_i <= '0';
                when 2095 => sda_i <= '0';
                when 2096 => sda_i <= '0';
                when 2097 => sda_i <= '0';
                when 2098 => sda_i <= '0';
                when 2099 => sda_i <= '0';
                when 2100 => sda_i <= '0';
                when 2101 => sda_i <= '0';
                when 2102 => sda_i <= '0';
                when 2103 => sda_i <= '0';
                when 2104 => sda_i <= '0';
                when 2105 => sda_i <= '0';
                when 2106 => sda_i <= '0';
                when 2107 => sda_i <= '0';
                when 2108 => sda_i <= '0';
                when 2109 => sda_i <= '0';
                when 2110 => sda_i <= '0';
                when 2111 => sda_i <= '0';
                when 2112 => sda_i <= '0';
                when 2113 => sda_i <= '0';
                when 2114 => sda_i <= '0';
                when 2115 => sda_i <= '0';
                when 2116 => sda_i <= '0';
                when 2117 => sda_i <= '0';
                when 2118 => sda_i <= '0';
                when 2119 => sda_i <= '0';
                when 2120 => sda_i <= '0';
                when 2121 => sda_i <= '0';
                when 2122 => sda_i <= '0';
                when 2123 => sda_i <= '0';
                when 2124 => sda_i <= '0';
                when 2125 => sda_i <= '0';
                when 2126 => sda_i <= '0';
                when 2127 => sda_i <= '0';
                when 2128 => sda_i <= '0';
                when 2129 => sda_i <= '0';
                when 2130 => sda_i <= '0';
                when 2131 => sda_i <= '0';
                when 2132 => sda_i <= '0';
                when 2133 => sda_i <= '0';
                when 2134 => sda_i <= '0';
                when 2135 => sda_i <= '0';
                when 2136 => sda_i <= '0';
                when 2137 => sda_i <= '0';
                when 2138 => sda_i <= '0';
                when 2139 => sda_i <= '0';
                when 2140 => sda_i <= '0';
                when 2141 => sda_i <= '0';
                when 2142 => sda_i <= '0';
                when 2143 => sda_i <= '0';
                when 2144 => sda_i <= '0';
                when 2145 => sda_i <= '0';
                when 2146 => sda_i <= '0';
                when 2147 => sda_i <= '0';
                when 2148 => sda_i <= '0';
                when 2149 => sda_i <= '0';
                when 2150 => sda_i <= '0';
                when 2151 => sda_i <= '0';
                when 2152 => sda_i <= '0';
                when 2153 => sda_i <= '0';
                when 2154 => sda_i <= '0';
                when 2155 => sda_i <= '0';
                when 2156 => sda_i <= '0';
                when 2157 => sda_i <= '0';
                when 2158 => sda_i <= '1';
                when 2159 => sda_i <= '1';
                when 2160 => sda_i <= '0';
                when 2161 => sda_i <= '0';
                when 2162 => sda_i <= '0';
                when 2163 => sda_i <= '0';
                when 2164 => sda_i <= '0';
                when 2165 => sda_i <= '0';
                when 2166 => sda_i <= '0';
                when 2167 => sda_i <= '0';
                when 2168 => sda_i <= '0';
                when 2169 => sda_i <= '0';
                when 2170 => sda_i <= '0';
                when 2171 => sda_i <= '0';
                when 2172 => sda_i <= '0';
                when 2173 => sda_i <= '0';
                when 2174 => sda_i <= '0';
                when 2175 => sda_i <= '0';
                when 2176 => sda_i <= '0';
                when 2177 => sda_i <= '0';
                when 2178 => sda_i <= '0';
                when 2179 => sda_i <= '0';
                when 2180 => sda_i <= '0';
                when 2181 => sda_i <= '0';
                when 2182 => sda_i <= '0';
                when 2183 => sda_i <= '0';
                when 2184 => sda_i <= '0';
                when 2185 => sda_i <= '0';
                when 2186 => sda_i <= '0';
                when 2187 => sda_i <= '0';
                when 2188 => sda_i <= '0';
                when 2189 => sda_i <= '0';
                when 2190 => sda_i <= '0';
                when 2191 => sda_i <= '0';
                when 2192 => sda_i <= '0';
                when 2193 => sda_i <= '0';
                when 2194 => sda_i <= '0';
                when 2195 => sda_i <= '0';
                when 2196 => sda_i <= '0';
                when 2197 => sda_i <= '0';
                when 2198 => sda_i <= '0';
                when 2199 => sda_i <= '0';
                when 2200 => sda_i <= '0';
                when 2201 => sda_i <= '0';
                when 2202 => sda_i <= '0';
                when 2203 => sda_i <= '0';
                when 2204 => sda_i <= '0';
                when 2205 => sda_i <= '0';
                when 2206 => sda_i <= '0';
                when 2207 => sda_i <= '0';
                when 2208 => sda_i <= '0';
                when 2209 => sda_i <= '0';
                when 2210 => sda_i <= '0';
                when 2211 => sda_i <= '0';
                when 2212 => sda_i <= '0';
                when 2213 => sda_i <= '0';
                when 2214 => sda_i <= '0';
                when 2215 => sda_i <= '0';
                when 2216 => sda_i <= '0';
                when 2217 => sda_i <= '0';
                when 2218 => sda_i <= '0';
                when 2219 => sda_i <= '0';
                when 2220 => sda_i <= '0';
                when 2221 => sda_i <= '0';
                when 2222 => sda_i <= '0';
                when 2223 => sda_i <= '0';
                when 2224 => sda_i <= '0';
                when 2225 => sda_i <= '0';
                when 2226 => sda_i <= '0';
                when 2227 => sda_i <= '0';
                when 2228 => sda_i <= '0';
                when 2229 => sda_i <= '0';
                when 2230 => sda_i <= '0';
                when 2231 => sda_i <= '0';
                when 2232 => sda_i <= '0';
                when 2233 => sda_i <= '0';
                when 2234 => sda_i <= '0';
                when 2235 => sda_i <= '0';
                when 2236 => sda_i <= '0';
                when 2237 => sda_i <= '0';
                when 2238 => sda_i <= '0';
                when 2239 => sda_i <= '0';
                when 2240 => sda_i <= '0';
                when 2241 => sda_i <= '0';
                when 2242 => sda_i <= '0';
                when 2243 => sda_i <= '0';
                when 2244 => sda_i <= '0';
                when 2245 => sda_i <= '0';
                when 2246 => sda_i <= '0';
                when 2247 => sda_i <= '0';
                when 2248 => sda_i <= '0';
                when 2249 => sda_i <= '0';
                when 2250 => sda_i <= '0';
                when 2251 => sda_i <= '0';
                when 2252 => sda_i <= '0';
                when 2253 => sda_i <= '0';
                when 2254 => sda_i <= '0';
                when 2255 => sda_i <= '0';
                when 2256 => sda_i <= '0';
                when 2257 => sda_i <= '0';
                when 2258 => sda_i <= '0';
                when 2259 => sda_i <= '0';
                when 2260 => sda_i <= '0';
                when 2261 => sda_i <= '0';
                when 2262 => sda_i <= '0';
                when 2263 => sda_i <= '0';
                when 2264 => sda_i <= '0';
                when 2265 => sda_i <= '0';
                when 2266 => sda_i <= '1';
                when 2267 => sda_i <= '1';
                when 2268 => sda_i <= '0';
                when 2269 => sda_i <= '0';
                when 2270 => sda_i <= '0';
                when 2271 => sda_i <= '0';
                when 2272 => sda_i <= '0';
                when 2273 => sda_i <= '0';
                when 2274 => sda_i <= '0';
                when 2275 => sda_i <= '0';
                when 2276 => sda_i <= '0';
                when 2277 => sda_i <= '0';
                when 2278 => sda_i <= '0';
                when 2279 => sda_i <= '0';
                when 2280 => sda_i <= '0';
                when 2281 => sda_i <= '0';
                when 2282 => sda_i <= '0';
                when 2283 => sda_i <= '0';
                when 2284 => sda_i <= '0';
                when 2285 => sda_i <= '0';
                when 2286 => sda_i <= '0';
                when 2287 => sda_i <= '0';
                when 2288 => sda_i <= '0';
                when 2289 => sda_i <= '0';
                when 2290 => sda_i <= '0';
                when 2291 => sda_i <= '0';
                when 2292 => sda_i <= '0';
                when 2293 => sda_i <= '0';
                when 2294 => sda_i <= '0';
                when 2295 => sda_i <= '0';
                when 2296 => sda_i <= '0';
                when 2297 => sda_i <= '0';
                when 2298 => sda_i <= '0';
                when 2299 => sda_i <= '0';
                when 2300 => sda_i <= '0';
                when 2301 => sda_i <= '0';
                when 2302 => sda_i <= '0';
                when 2303 => sda_i <= '0';
                when 2304 => sda_i <= '0';
                when 2305 => sda_i <= '0';
                when 2306 => sda_i <= '0';
                when 2307 => sda_i <= '0';
                when 2308 => sda_i <= '0';
                when 2309 => sda_i <= '0';
                when 2310 => sda_i <= '0';
                when 2311 => sda_i <= '0';
                when 2312 => sda_i <= '0';
                when 2313 => sda_i <= '0';
                when 2314 => sda_i <= '0';
                when 2315 => sda_i <= '0';
                when 2316 => sda_i <= '0';
                when 2317 => sda_i <= '0';
                when 2318 => sda_i <= '0';
                when 2319 => sda_i <= '0';
                when 2320 => sda_i <= '0';
                when 2321 => sda_i <= '0';
                when 2322 => sda_i <= '0';
                when 2323 => sda_i <= '0';
                when 2324 => sda_i <= '0';
                when 2325 => sda_i <= '0';
                when 2326 => sda_i <= '0';
                when 2327 => sda_i <= '0';
                when 2328 => sda_i <= '0';
                when 2329 => sda_i <= '0';
                when 2330 => sda_i <= '0';
                when 2331 => sda_i <= '0';
                when 2332 => sda_i <= '0';
                when 2333 => sda_i <= '0';
                when 2334 => sda_i <= '0';
                when 2335 => sda_i <= '0';
                when 2336 => sda_i <= '0';
                when 2337 => sda_i <= '0';
                when 2338 => sda_i <= '0';
                when 2339 => sda_i <= '0';
                when 2340 => sda_i <= '0';
                when 2341 => sda_i <= '0';
                when 2342 => sda_i <= '0';
                when 2343 => sda_i <= '0';
                when 2344 => sda_i <= '0';
                when 2345 => sda_i <= '0';
                when 2346 => sda_i <= '0';
                when 2347 => sda_i <= '0';
                when 2348 => sda_i <= '0';
                when 2349 => sda_i <= '0';
                when 2350 => sda_i <= '0';
                when 2351 => sda_i <= '0';
                when 2352 => sda_i <= '0';
                when 2353 => sda_i <= '0';
                when 2354 => sda_i <= '0';
                when 2355 => sda_i <= '0';
                when 2356 => sda_i <= '0';
                when 2357 => sda_i <= '0';
                when 2358 => sda_i <= '0';
                when 2359 => sda_i <= '0';
                when 2360 => sda_i <= '0';
                when 2361 => sda_i <= '0';
                when 2362 => sda_i <= '0';
                when 2363 => sda_i <= '0';
                when 2364 => sda_i <= '0';
                when 2365 => sda_i <= '0';
                when 2366 => sda_i <= '0';
                when 2367 => sda_i <= '0';
                when 2368 => sda_i <= '0';
                when 2369 => sda_i <= '0';
                when 2370 => sda_i <= '0';
                when 2371 => sda_i <= '0';
                when 2372 => sda_i <= '0';
                when 2373 => sda_i <= '0';
                when 2374 => sda_i <= '1';
                when 2375 => sda_i <= '1';
                when 2376 => sda_i <= '0';
                when 2377 => sda_i <= '0';
                when 2378 => sda_i <= '0';
                when 2379 => sda_i <= '0';
                when 2380 => sda_i <= '0';
                when 2381 => sda_i <= '0';
                when 2382 => sda_i <= '0';
                when 2383 => sda_i <= '0';
                when 2384 => sda_i <= '0';
                when 2385 => sda_i <= '0';
                when 2386 => sda_i <= '0';
                when 2387 => sda_i <= '0';
                when 2388 => sda_i <= '0';
                when 2389 => sda_i <= '0';
                when 2390 => sda_i <= '0';
                when 2391 => sda_i <= '0';
                when 2392 => sda_i <= '0';
                when 2393 => sda_i <= '0';
                when 2394 => sda_i <= '0';
                when 2395 => sda_i <= '0';
                when 2396 => sda_i <= '0';
                when 2397 => sda_i <= '0';
                when 2398 => sda_i <= '0';
                when 2399 => sda_i <= '0';
                when 2400 => sda_i <= '0';
                when 2401 => sda_i <= '0';
                when 2402 => sda_i <= '0';
                when 2403 => sda_i <= '0';
                when 2404 => sda_i <= '0';
                when 2405 => sda_i <= '0';
                when 2406 => sda_i <= '0';
                when 2407 => sda_i <= '0';
                when 2408 => sda_i <= '0';
                when 2409 => sda_i <= '0';
                when 2410 => sda_i <= '0';
                when 2411 => sda_i <= '0';
                when 2412 => sda_i <= '0';
                when 2413 => sda_i <= '0';
                when 2414 => sda_i <= '0';
                when 2415 => sda_i <= '0';
                when 2416 => sda_i <= '0';
                when 2417 => sda_i <= '0';
                when 2418 => sda_i <= '0';
                when 2419 => sda_i <= '0';
                when 2420 => sda_i <= '0';
                when 2421 => sda_i <= '0';
                when 2422 => sda_i <= '0';
                when 2423 => sda_i <= '0';
                when 2424 => sda_i <= '0';
                when 2425 => sda_i <= '0';
                when 2426 => sda_i <= '0';
                when 2427 => sda_i <= '0';
                when 2428 => sda_i <= '0';
                when 2429 => sda_i <= '0';
                when 2430 => sda_i <= '0';
                when 2431 => sda_i <= '0';
                when 2432 => sda_i <= '0';
                when 2433 => sda_i <= '0';
                when 2434 => sda_i <= '0';
                when 2435 => sda_i <= '0';
                when 2436 => sda_i <= '0';
                when 2437 => sda_i <= '0';
                when 2438 => sda_i <= '0';
                when 2439 => sda_i <= '0';
                when 2440 => sda_i <= '0';
                when 2441 => sda_i <= '0';
                when 2442 => sda_i <= '0';
                when 2443 => sda_i <= '0';
                when 2444 => sda_i <= '0';
                when 2445 => sda_i <= '0';
                when 2446 => sda_i <= '0';
                when 2447 => sda_i <= '0';
                when 2448 => sda_i <= '0';
                when 2449 => sda_i <= '0';
                when 2450 => sda_i <= '0';
                when 2451 => sda_i <= '0';
                when 2452 => sda_i <= '0';
                when 2453 => sda_i <= '0';
                when 2454 => sda_i <= '0';
                when 2455 => sda_i <= '0';
                when 2456 => sda_i <= '0';
                when 2457 => sda_i <= '0';
                when 2458 => sda_i <= '0';
                when 2459 => sda_i <= '0';
                when 2460 => sda_i <= '0';
                when 2461 => sda_i <= '0';
                when 2462 => sda_i <= '0';
                when 2463 => sda_i <= '0';
                when 2464 => sda_i <= '0';
                when 2465 => sda_i <= '0';
                when 2466 => sda_i <= '0';
                when 2467 => sda_i <= '0';
                when 2468 => sda_i <= '0';
                when 2469 => sda_i <= '0';
                when 2470 => sda_i <= '0';
                when 2471 => sda_i <= '0';
                when 2472 => sda_i <= '0';
                when 2473 => sda_i <= '0';
                when 2474 => sda_i <= '0';
                when 2475 => sda_i <= '0';
                when 2476 => sda_i <= '0';
                when 2477 => sda_i <= '0';
                when 2478 => sda_i <= '0';
                when 2479 => sda_i <= '0';
                when 2480 => sda_i <= '0';
                when 2481 => sda_i <= '0';
                when 2482 => sda_i <= '1';
                when 2483 => sda_i <= '1';
                when 2484 => sda_i <= '0';
                when 2485 => sda_i <= '0';
                when 2486 => sda_i <= '0';
                when 2487 => sda_i <= '0';
                when 2488 => sda_i <= '0';
                when 2489 => sda_i <= '0';
                when 2490 => sda_i <= '0';
                when 2491 => sda_i <= '0';
                when 2492 => sda_i <= '0';
                when 2493 => sda_i <= '0';
                when 2494 => sda_i <= '0';
                when 2495 => sda_i <= '0';
                when 2496 => sda_i <= '0';
                when 2497 => sda_i <= '0';
                when 2498 => sda_i <= '0';
                when 2499 => sda_i <= '0';
                when 2500 => sda_i <= '0';
                when 2501 => sda_i <= '0';
                when 2502 => sda_i <= '0';
                when 2503 => sda_i <= '0';
                when 2504 => sda_i <= '0';
                when 2505 => sda_i <= '0';
                when 2506 => sda_i <= '0';
                when 2507 => sda_i <= '0';
                when 2508 => sda_i <= '0';
                when 2509 => sda_i <= '0';
                when 2510 => sda_i <= '0';
                when 2511 => sda_i <= '0';
                when 2512 => sda_i <= '0';
                when 2513 => sda_i <= '0';
                when 2514 => sda_i <= '0';
                when 2515 => sda_i <= '0';
                when 2516 => sda_i <= '0';
                when 2517 => sda_i <= '0';
                when 2518 => sda_i <= '0';
                when 2519 => sda_i <= '0';
                when 2520 => sda_i <= '0';
                when 2521 => sda_i <= '0';
                when 2522 => sda_i <= '0';
                when 2523 => sda_i <= '0';
                when 2524 => sda_i <= '0';
                when 2525 => sda_i <= '0';
                when 2526 => sda_i <= '0';
                when 2527 => sda_i <= '0';
                when 2528 => sda_i <= '0';
                when 2529 => sda_i <= '0';
                when 2530 => sda_i <= '0';
                when 2531 => sda_i <= '0';
                when 2532 => sda_i <= '0';
                when 2533 => sda_i <= '0';
                when 2534 => sda_i <= '0';
                when 2535 => sda_i <= '0';
                when 2536 => sda_i <= '0';
                when 2537 => sda_i <= '0';
                when 2538 => sda_i <= '0';
                when 2539 => sda_i <= '0';
                when 2540 => sda_i <= '0';
                when 2541 => sda_i <= '0';
                when 2542 => sda_i <= '0';
                when 2543 => sda_i <= '0';
                when 2544 => sda_i <= '0';
                when 2545 => sda_i <= '0';
                when 2546 => sda_i <= '0';
                when 2547 => sda_i <= '0';
                when 2548 => sda_i <= '0';
                when 2549 => sda_i <= '0';
                when 2550 => sda_i <= '0';
                when 2551 => sda_i <= '0';
                when 2552 => sda_i <= '0';
                when 2553 => sda_i <= '0';
                when 2554 => sda_i <= '0';
                when 2555 => sda_i <= '0';
                when 2556 => sda_i <= '0';
                when 2557 => sda_i <= '0';
                when 2558 => sda_i <= '0';
                when 2559 => sda_i <= '0';
                when 2560 => sda_i <= '0';
                when 2561 => sda_i <= '0';
                when 2562 => sda_i <= '0';
                when 2563 => sda_i <= '0';
                when 2564 => sda_i <= '0';
                when 2565 => sda_i <= '0';
                when 2566 => sda_i <= '0';
                when 2567 => sda_i <= '0';
                when 2568 => sda_i <= '0';
                when 2569 => sda_i <= '0';
                when 2570 => sda_i <= '0';
                when 2571 => sda_i <= '0';
                when 2572 => sda_i <= '0';
                when 2573 => sda_i <= '0';
                when 2574 => sda_i <= '0';
                when 2575 => sda_i <= '0';
                when 2576 => sda_i <= '0';
                when 2577 => sda_i <= '0';
                when 2578 => sda_i <= '0';
                when 2579 => sda_i <= '0';
                when 2580 => sda_i <= '0';
                when 2581 => sda_i <= '0';
                when 2582 => sda_i <= '0';
                when 2583 => sda_i <= '0';
                when 2584 => sda_i <= '0';
                when 2585 => sda_i <= '0';
                when 2586 => sda_i <= '0';
                when 2587 => sda_i <= '0';
                when 2588 => sda_i <= '0';
                when 2589 => sda_i <= '0';
                when 2590 => sda_i <= '1';
                when 2591 => sda_i <= '1';
                when 2592 => sda_i <= '0';
                when 2593 => sda_i <= '0';
                when 2594 => sda_i <= '0';
                when 2595 => sda_i <= '0';
                when 2596 => sda_i <= '0';
                when 2597 => sda_i <= '0';
                when 2598 => sda_i <= '0';
                when 2599 => sda_i <= '0';
                when 2600 => sda_i <= '0';
                when 2601 => sda_i <= '0';
                when 2602 => sda_i <= '0';
                when 2603 => sda_i <= '0';
                when 2604 => sda_i <= '0';
                when 2605 => sda_i <= '0';
                when 2606 => sda_i <= '0';
                when 2607 => sda_i <= '0';
                when 2608 => sda_i <= '0';
                when 2609 => sda_i <= '0';
                when 2610 => sda_i <= '0';
                when 2611 => sda_i <= '0';
                when 2612 => sda_i <= '0';
                when 2613 => sda_i <= '0';
                when 2614 => sda_i <= '0';
                when 2615 => sda_i <= '0';
                when 2616 => sda_i <= '0';
                when 2617 => sda_i <= '0';
                when 2618 => sda_i <= '0';
                when 2619 => sda_i <= '0';
                when 2620 => sda_i <= '0';
                when 2621 => sda_i <= '0';
                when 2622 => sda_i <= '0';
                when 2623 => sda_i <= '0';
                when 2624 => sda_i <= '0';
                when 2625 => sda_i <= '0';
                when 2626 => sda_i <= '0';
                when 2627 => sda_i <= '0';
                when 2628 => sda_i <= '0';
                when 2629 => sda_i <= '0';
                when 2630 => sda_i <= '0';
                when 2631 => sda_i <= '0';
                when 2632 => sda_i <= '0';
                when 2633 => sda_i <= '0';
                when 2634 => sda_i <= '0';
                when 2635 => sda_i <= '0';
                when 2636 => sda_i <= '0';
                when 2637 => sda_i <= '0';
                when 2638 => sda_i <= '0';
                when 2639 => sda_i <= '0';
                when 2640 => sda_i <= '0';
                when 2641 => sda_i <= '0';
                when 2642 => sda_i <= '0';
                when 2643 => sda_i <= '0';
                when 2644 => sda_i <= '0';
                when 2645 => sda_i <= '0';
                when 2646 => sda_i <= '0';
                when 2647 => sda_i <= '0';
                when 2648 => sda_i <= '0';
                when 2649 => sda_i <= '0';
                when 2650 => sda_i <= '0';
                when 2651 => sda_i <= '0';
                when 2652 => sda_i <= '0';
                when 2653 => sda_i <= '0';
                when 2654 => sda_i <= '0';
                when 2655 => sda_i <= '0';
                when 2656 => sda_i <= '0';
                when 2657 => sda_i <= '0';
                when 2658 => sda_i <= '0';
                when 2659 => sda_i <= '0';
                when 2660 => sda_i <= '0';
                when 2661 => sda_i <= '0';
                when 2662 => sda_i <= '0';
                when 2663 => sda_i <= '0';
                when 2664 => sda_i <= '0';
                when 2665 => sda_i <= '0';
                when 2666 => sda_i <= '0';
                when 2667 => sda_i <= '0';
                when 2668 => sda_i <= '0';
                when 2669 => sda_i <= '0';
                when 2670 => sda_i <= '0';
                when 2671 => sda_i <= '0';
                when 2672 => sda_i <= '0';
                when 2673 => sda_i <= '0';
                when 2674 => sda_i <= '0';
                when 2675 => sda_i <= '0';
                when 2676 => sda_i <= '0';
                when 2677 => sda_i <= '0';
                when 2678 => sda_i <= '0';
                when 2679 => sda_i <= '0';
                when 2680 => sda_i <= '0';
                when 2681 => sda_i <= '0';
                when 2682 => sda_i <= '0';
                when 2683 => sda_i <= '0';
                when 2684 => sda_i <= '0';
                when 2685 => sda_i <= '0';
                when 2686 => sda_i <= '0';
                when 2687 => sda_i <= '0';
                when 2688 => sda_i <= '0';
                when 2689 => sda_i <= '0';
                when 2690 => sda_i <= '0';
                when 2691 => sda_i <= '0';
                when 2692 => sda_i <= '0';
                when 2693 => sda_i <= '0';
                when 2694 => sda_i <= '0';
                when 2695 => sda_i <= '0';
                when 2696 => sda_i <= '0';
                when 2697 => sda_i <= '0';
                when 2698 => sda_i <= '1';
                when 2699 => sda_i <= '1';
                when 2700 => sda_i <= '0';
                when 2701 => sda_i <= '0';
                when 2702 => sda_i <= '0';
                when 2703 => sda_i <= '0';
                when 2704 => sda_i <= '0';
                when 2705 => sda_i <= '0';
                when 2706 => sda_i <= '0';
                when 2707 => sda_i <= '0';
                when 2708 => sda_i <= '0';
                when 2709 => sda_i <= '0';
                when 2710 => sda_i <= '0';
                when 2711 => sda_i <= '0';
                when 2712 => sda_i <= '0';
                when 2713 => sda_i <= '0';
                when 2714 => sda_i <= '0';
                when 2715 => sda_i <= '0';
                when 2716 => sda_i <= '0';
                when 2717 => sda_i <= '0';
                when 2718 => sda_i <= '0';
                when 2719 => sda_i <= '0';
                when 2720 => sda_i <= '0';
                when 2721 => sda_i <= '0';
                when 2722 => sda_i <= '0';
                when 2723 => sda_i <= '0';
                when 2724 => sda_i <= '0';
                when 2725 => sda_i <= '0';
                when 2726 => sda_i <= '0';
                when 2727 => sda_i <= '0';
                when 2728 => sda_i <= '0';
                when 2729 => sda_i <= '0';
                when 2730 => sda_i <= '0';
                when 2731 => sda_i <= '0';
                when 2732 => sda_i <= '0';
                when 2733 => sda_i <= '0';
                when 2734 => sda_i <= '0';
                when 2735 => sda_i <= '0';
                when 2736 => sda_i <= '0';
                when 2737 => sda_i <= '0';
                when 2738 => sda_i <= '0';
                when 2739 => sda_i <= '0';
                when 2740 => sda_i <= '0';
                when 2741 => sda_i <= '0';
                when 2742 => sda_i <= '0';
                when 2743 => sda_i <= '0';
                when 2744 => sda_i <= '0';
                when 2745 => sda_i <= '0';
                when 2746 => sda_i <= '0';
                when 2747 => sda_i <= '0';
                when 2748 => sda_i <= '0';
                when 2749 => sda_i <= '0';
                when 2750 => sda_i <= '0';
                when 2751 => sda_i <= '0';
                when 2752 => sda_i <= '0';
                when 2753 => sda_i <= '0';
                when 2754 => sda_i <= '0';
                when 2755 => sda_i <= '0';
                when 2756 => sda_i <= '0';
                when 2757 => sda_i <= '0';
                when 2758 => sda_i <= '0';
                when 2759 => sda_i <= '0';
                when 2760 => sda_i <= '0';
                when 2761 => sda_i <= '0';
                when 2762 => sda_i <= '0';
                when 2763 => sda_i <= '0';
                when 2764 => sda_i <= '0';
                when 2765 => sda_i <= '0';
                when 2766 => sda_i <= '0';
                when 2767 => sda_i <= '0';
                when 2768 => sda_i <= '0';
                when 2769 => sda_i <= '0';
                when 2770 => sda_i <= '0';
                when 2771 => sda_i <= '0';
                when 2772 => sda_i <= '0';
                when 2773 => sda_i <= '0';
                when 2774 => sda_i <= '0';
                when 2775 => sda_i <= '0';
                when 2776 => sda_i <= '0';
                when 2777 => sda_i <= '0';
                when 2778 => sda_i <= '0';
                when 2779 => sda_i <= '0';
                when 2780 => sda_i <= '0';
                when 2781 => sda_i <= '0';
                when 2782 => sda_i <= '0';
                when 2783 => sda_i <= '0';
                when 2784 => sda_i <= '0';
                when 2785 => sda_i <= '0';
                when 2786 => sda_i <= '0';
                when 2787 => sda_i <= '0';
                when 2788 => sda_i <= '0';
                when 2789 => sda_i <= '0';
                when 2790 => sda_i <= '0';
                when 2791 => sda_i <= '0';
                when 2792 => sda_i <= '0';
                when 2793 => sda_i <= '0';
                when 2794 => sda_i <= '0';
                when 2795 => sda_i <= '0';
                when 2796 => sda_i <= '0';
                when 2797 => sda_i <= '0';
                when 2798 => sda_i <= '0';
                when 2799 => sda_i <= '0';
                when 2800 => sda_i <= '0';
                when 2801 => sda_i <= '0';
                when 2802 => sda_i <= '0';
                when 2803 => sda_i <= '0';
                when 2804 => sda_i <= '0';
                when 2805 => sda_i <= '0';
                when 2806 => sda_i <= '1';
                when 2807 => sda_i <= '1';
                when 2808 => sda_i <= '0';
                when 2809 => sda_i <= '0';
                when 2810 => sda_i <= '0';
                when 2811 => sda_i <= '0';
                when 2812 => sda_i <= '0';
                when 2813 => sda_i <= '0';
                when 2814 => sda_i <= '0';
                when 2815 => sda_i <= '0';
                when 2816 => sda_i <= '0';
                when 2817 => sda_i <= '0';
                when 2818 => sda_i <= '0';
                when 2819 => sda_i <= '0';
                when 2820 => sda_i <= '1';
                when 2821 => sda_i <= '1';
                when 2822 => sda_i <= '1';
                when 2823 => sda_i <= '1';
                when 2824 => sda_i <= '1';
                when 2825 => sda_i <= '1';
                when 2826 => sda_i <= '1';
                when 2827 => sda_i <= '1';
                when 2828 => sda_i <= '1';
                when 2829 => sda_i <= '1';
                when 2830 => sda_i <= '1';
                when 2831 => sda_i <= '1';
                when 2832 => sda_i <= '1';
                when 2833 => sda_i <= '1';
                when 2834 => sda_i <= '1';
                when 2835 => sda_i <= '1';
                when 2836 => sda_i <= '1';
                when 2837 => sda_i <= '1';
                when 2838 => sda_i <= '1';
                when 2839 => sda_i <= '1';
                when 2840 => sda_i <= '1';
                when 2841 => sda_i <= '1';
                when 2842 => sda_i <= '1';
                when 2843 => sda_i <= '1';
                when 2844 => sda_i <= '1';
                when 2845 => sda_i <= '1';
                when 2846 => sda_i <= '1';
                when 2847 => sda_i <= '1';
                when 2848 => sda_i <= '1';
                when 2849 => sda_i <= '1';
                when 2850 => sda_i <= '1';
                when 2851 => sda_i <= '1';
                when 2852 => sda_i <= '1';
                when 2853 => sda_i <= '0';
                when 2854 => sda_i <= '0';
                when 2855 => sda_i <= '0';
                when 2856 => sda_i <= '0';
                when 2857 => sda_i <= '0';
                when 2858 => sda_i <= '0';
                when 2859 => sda_i <= '0';
                when 2860 => sda_i <= '0';
                when 2861 => sda_i <= '0';
                when 2862 => sda_i <= '0';
                when 2863 => sda_i <= '0';
                when 2864 => sda_i <= '0';
                when 2865 => sda_i <= '0';
                when 2866 => sda_i <= '0';
                when 2867 => sda_i <= '0';
                when 2868 => sda_i <= '0';
                when 2869 => sda_i <= '0';
                when 2870 => sda_i <= '0';
                when 2871 => sda_i <= '0';
                when 2872 => sda_i <= '0';
                when 2873 => sda_i <= '0';
                when 2874 => sda_i <= '0';
                when 2875 => sda_i <= '0';
                when 2876 => sda_i <= '0';
                when 2877 => sda_i <= '0';
                when 2878 => sda_i <= '1';
                when 2879 => sda_i <= '1';
                when 2880 => sda_i <= '1';
                when 2881 => sda_i <= '1';
                when 2882 => sda_i <= '1';
                when 2883 => sda_i <= '1';
                when 2884 => sda_i <= '1';
                when 2885 => sda_i <= '1';
                when 2886 => sda_i <= '1';
                when 2887 => sda_i <= '1';
                when 2888 => sda_i <= '1';
                when 2889 => sda_i <= '0';
                when 2890 => sda_i <= '0';
                when 2891 => sda_i <= '0';
                when 2892 => sda_i <= '0';
                when 2893 => sda_i <= '0';
                when 2894 => sda_i <= '0';
                when 2895 => sda_i <= '0';
                when 2896 => sda_i <= '0';
                when 2897 => sda_i <= '0';
                when 2898 => sda_i <= '0';
                when 2899 => sda_i <= '0';
                when 2900 => sda_i <= '0';
                when 2901 => sda_i <= '0';
                when 2902 => sda_i <= '1';
                when 2903 => sda_i <= '1';
                when 2904 => sda_i <= '1';
                when 2905 => sda_i <= '1';
                when 2906 => sda_i <= '1';
                when 2907 => sda_i <= '1';
                when 2908 => sda_i <= '1';
                when 2909 => sda_i <= '1';
                when 2910 => sda_i <= '1';
                when 2911 => sda_i <= '1';
                when 2912 => sda_i <= '1';
                when 2913 => sda_i <= '1';
                when 2914 => sda_i <= '1';
                when 2915 => sda_i <= '1';
                when 2916 => sda_i <= '0';
                when 2917 => sda_i <= '0';
                when 2918 => sda_i <= '0';
                when 2919 => sda_i <= '0';
                when 2920 => sda_i <= '0';
                when 2921 => sda_i <= '0';
                when 2922 => sda_i <= '0';
                when 2923 => sda_i <= '0';
                when 2924 => sda_i <= '0';
                when 2925 => sda_i <= '0';
                when 2926 => sda_i <= '0';
                when 2927 => sda_i <= '0';
                when 2928 => sda_i <= '0';
                when 2929 => sda_i <= '0';
                when 2930 => sda_i <= '0';
                when 2931 => sda_i <= '0';
                when 2932 => sda_i <= '0';
                when 2933 => sda_i <= '0';
                when 2934 => sda_i <= '0';
                when 2935 => sda_i <= '0';
                when 2936 => sda_i <= '0';
                when 2937 => sda_i <= '0';
                when 2938 => sda_i <= '0';
                when 2939 => sda_i <= '0';
                when 2940 => sda_i <= '0';
                when 2941 => sda_i <= '0';
                when 2942 => sda_i <= '0';
                when 2943 => sda_i <= '0';
                when 2944 => sda_i <= '0';
                when 2945 => sda_i <= '0';
                when 2946 => sda_i <= '0';
                when 2947 => sda_i <= '0';
                when 2948 => sda_i <= '0';
                when 2949 => sda_i <= '0';
                when 2950 => sda_i <= '0';
                when 2951 => sda_i <= '0';
                when 2952 => sda_i <= '0';
                when 2953 => sda_i <= '0';
                when 2954 => sda_i <= '0';
                when 2955 => sda_i <= '0';
                when 2956 => sda_i <= '0';
                when 2957 => sda_i <= '0';
                when 2958 => sda_i <= '0';
                when 2959 => sda_i <= '0';
                when 2960 => sda_i <= '0';
                when 2961 => sda_i <= '0';
                when 2962 => sda_i <= '0';
                when 2963 => sda_i <= '0';
                when 2964 => sda_i <= '0';
                when 2965 => sda_i <= '0';
                when 2966 => sda_i <= '0';
                when 2967 => sda_i <= '0';
                when 2968 => sda_i <= '0';
                when 2969 => sda_i <= '0';
                when 2970 => sda_i <= '0';
                when 2971 => sda_i <= '0';
                when 2972 => sda_i <= '0';
                when 2973 => sda_i <= '0';
                when 2974 => sda_i <= '0';
                when 2975 => sda_i <= '0';
                when 2976 => sda_i <= '0';
                when 2977 => sda_i <= '0';
                when 2978 => sda_i <= '0';
                when 2979 => sda_i <= '0';
                when 2980 => sda_i <= '0';
                when 2981 => sda_i <= '0';
                when 2982 => sda_i <= '0';
                when 2983 => sda_i <= '0';
                when 2984 => sda_i <= '0';
                when 2985 => sda_i <= '0';
                when 2986 => sda_i <= '0';
                when 2987 => sda_i <= '0';
                when 2988 => sda_i <= '0';
                when 2989 => sda_i <= '0';
                when 2990 => sda_i <= '0';
                when 2991 => sda_i <= '0';
                when 2992 => sda_i <= '0';
                when 2993 => sda_i <= '0';
                when 2994 => sda_i <= '0';
                when 2995 => sda_i <= '0';
                when 2996 => sda_i <= '0';
                when 2997 => sda_i <= '0';
                when 2998 => sda_i <= '0';
                when 2999 => sda_i <= '0';
                when 3000 => sda_i <= '0';
                when 3001 => sda_i <= '0';
                when 3002 => sda_i <= '0';
                when 3003 => sda_i <= '0';
                when 3004 => sda_i <= '0';
                when 3005 => sda_i <= '0';
                when 3006 => sda_i <= '0';
                when 3007 => sda_i <= '0';
                when 3008 => sda_i <= '0';
                when 3009 => sda_i <= '0';
                when 3010 => sda_i <= '0';
                when 3011 => sda_i <= '0';
                when 3012 => sda_i <= '0';
                when 3013 => sda_i <= '0';
                when 3014 => sda_i <= '0';
                when 3015 => sda_i <= '0';
                when 3016 => sda_i <= '0';
                when 3017 => sda_i <= '0';
                when 3018 => sda_i <= '0';
                when 3019 => sda_i <= '0';
                when 3020 => sda_i <= '0';
                when 3021 => sda_i <= '0';
                when 3022 => sda_i <= '1';
                when 3023 => sda_i <= '1';
                when 3024 => sda_i <= '0';
                when 3025 => sda_i <= '0';
                when 3026 => sda_i <= '0';
                when 3027 => sda_i <= '0';
                when 3028 => sda_i <= '0';
                when 3029 => sda_i <= '0';
                when 3030 => sda_i <= '0';
                when 3031 => sda_i <= '0';
                when 3032 => sda_i <= '0';
                when 3033 => sda_i <= '0';
                when 3034 => sda_i <= '0';
                when 3035 => sda_i <= '0';
                when 3036 => sda_i <= '0';
                when 3037 => sda_i <= '0';
                when 3038 => sda_i <= '0';
                when 3039 => sda_i <= '0';
                when 3040 => sda_i <= '0';
                when 3041 => sda_i <= '0';
                when 3042 => sda_i <= '0';
                when 3043 => sda_i <= '0';
                when 3044 => sda_i <= '0';
                when 3045 => sda_i <= '0';
                when 3046 => sda_i <= '0';
                when 3047 => sda_i <= '0';
                when 3048 => sda_i <= '0';
                when 3049 => sda_i <= '0';
                when 3050 => sda_i <= '0';
                when 3051 => sda_i <= '0';
                when 3052 => sda_i <= '0';
                when 3053 => sda_i <= '0';
                when 3054 => sda_i <= '0';
                when 3055 => sda_i <= '0';
                when 3056 => sda_i <= '0';
                when 3057 => sda_i <= '0';
                when 3058 => sda_i <= '0';
                when 3059 => sda_i <= '0';
                when 3060 => sda_i <= '0';
                when 3061 => sda_i <= '0';
                when 3062 => sda_i <= '0';
                when 3063 => sda_i <= '0';
                when 3064 => sda_i <= '0';
                when 3065 => sda_i <= '0';
                when 3066 => sda_i <= '0';
                when 3067 => sda_i <= '0';
                when 3068 => sda_i <= '0';
                when 3069 => sda_i <= '0';
                when 3070 => sda_i <= '0';
                when 3071 => sda_i <= '0';
                when 3072 => sda_i <= '0';
                when 3073 => sda_i <= '0';
                when 3074 => sda_i <= '0';
                when 3075 => sda_i <= '0';
                when 3076 => sda_i <= '0';
                when 3077 => sda_i <= '0';
                when 3078 => sda_i <= '0';
                when 3079 => sda_i <= '0';
                when 3080 => sda_i <= '0';
                when 3081 => sda_i <= '0';
                when 3082 => sda_i <= '0';
                when 3083 => sda_i <= '0';
                when 3084 => sda_i <= '0';
                when 3085 => sda_i <= '0';
                when 3086 => sda_i <= '0';
                when 3087 => sda_i <= '0';
                when 3088 => sda_i <= '0';
                when 3089 => sda_i <= '0';
                when 3090 => sda_i <= '0';
                when 3091 => sda_i <= '0';
                when 3092 => sda_i <= '0';
                when 3093 => sda_i <= '0';
                when 3094 => sda_i <= '0';
                when 3095 => sda_i <= '0';
                when 3096 => sda_i <= '0';
                when 3097 => sda_i <= '0';
                when 3098 => sda_i <= '0';
                when 3099 => sda_i <= '0';
                when 3100 => sda_i <= '0';
                when 3101 => sda_i <= '0';
                when 3102 => sda_i <= '0';
                when 3103 => sda_i <= '0';
                when 3104 => sda_i <= '0';
                when 3105 => sda_i <= '0';
                when 3106 => sda_i <= '0';
                when 3107 => sda_i <= '0';
                when 3108 => sda_i <= '0';
                when 3109 => sda_i <= '0';
                when 3110 => sda_i <= '0';
                when 3111 => sda_i <= '0';
                when 3112 => sda_i <= '0';
                when 3113 => sda_i <= '0';
                when 3114 => sda_i <= '0';
                when 3115 => sda_i <= '0';
                when 3116 => sda_i <= '0';
                when 3117 => sda_i <= '0';
                when 3118 => sda_i <= '0';
                when 3119 => sda_i <= '0';
                when 3120 => sda_i <= '0';
                when 3121 => sda_i <= '0';
                when 3122 => sda_i <= '0';
                when 3123 => sda_i <= '0';
                when 3124 => sda_i <= '0';
                when 3125 => sda_i <= '0';
                when 3126 => sda_i <= '0';
                when 3127 => sda_i <= '0';
                when 3128 => sda_i <= '0';
                when 3129 => sda_i <= '0';
                when 3130 => sda_i <= '1';
                when 3131 => sda_i <= '1';
                when 3132 => sda_i <= '0';
                when 3133 => sda_i <= '0';
                when 3134 => sda_i <= '0';
                when 3135 => sda_i <= '0';
                when 3136 => sda_i <= '0';
                when 3137 => sda_i <= '0';
                when 3138 => sda_i <= '0';
                when 3139 => sda_i <= '0';
                when 3140 => sda_i <= '0';
                when 3141 => sda_i <= '0';
                when 3142 => sda_i <= '0';
                when 3143 => sda_i <= '0';
                when 3144 => sda_i <= '0';
                when 3145 => sda_i <= '0';
                when 3146 => sda_i <= '0';
                when 3147 => sda_i <= '0';
                when 3148 => sda_i <= '0';
                when 3149 => sda_i <= '0';
                when 3150 => sda_i <= '0';
                when 3151 => sda_i <= '0';
                when 3152 => sda_i <= '0';
                when 3153 => sda_i <= '0';
                when 3154 => sda_i <= '0';
                when 3155 => sda_i <= '0';
                when 3156 => sda_i <= '0';
                when 3157 => sda_i <= '0';
                when 3158 => sda_i <= '0';
                when 3159 => sda_i <= '0';
                when 3160 => sda_i <= '0';
                when 3161 => sda_i <= '0';
                when 3162 => sda_i <= '0';
                when 3163 => sda_i <= '0';
                when 3164 => sda_i <= '0';
                when 3165 => sda_i <= '0';
                when 3166 => sda_i <= '0';
                when 3167 => sda_i <= '0';
                when 3168 => sda_i <= '0';
                when 3169 => sda_i <= '0';
                when 3170 => sda_i <= '0';
                when 3171 => sda_i <= '0';
                when 3172 => sda_i <= '0';
                when 3173 => sda_i <= '0';
                when 3174 => sda_i <= '0';
                when 3175 => sda_i <= '0';
                when 3176 => sda_i <= '0';
                when 3177 => sda_i <= '0';
                when 3178 => sda_i <= '0';
                when 3179 => sda_i <= '0';
                when 3180 => sda_i <= '0';
                when 3181 => sda_i <= '0';
                when 3182 => sda_i <= '0';
                when 3183 => sda_i <= '0';
                when 3184 => sda_i <= '0';
                when 3185 => sda_i <= '0';
                when 3186 => sda_i <= '0';
                when 3187 => sda_i <= '0';
                when 3188 => sda_i <= '0';
                when 3189 => sda_i <= '0';
                when 3190 => sda_i <= '0';
                when 3191 => sda_i <= '0';
                when 3192 => sda_i <= '0';
                when 3193 => sda_i <= '0';
                when 3194 => sda_i <= '0';
                when 3195 => sda_i <= '0';
                when 3196 => sda_i <= '0';
                when 3197 => sda_i <= '0';
                when 3198 => sda_i <= '0';
                when 3199 => sda_i <= '0';
                when 3200 => sda_i <= '0';
                when 3201 => sda_i <= '0';
                when 3202 => sda_i <= '0';
                when 3203 => sda_i <= '0';
                when 3204 => sda_i <= '0';
                when 3205 => sda_i <= '0';
                when 3206 => sda_i <= '0';
                when 3207 => sda_i <= '0';
                when 3208 => sda_i <= '0';
                when 3209 => sda_i <= '0';
                when 3210 => sda_i <= '0';
                when 3211 => sda_i <= '0';
                when 3212 => sda_i <= '0';
                when 3213 => sda_i <= '0';
                when 3214 => sda_i <= '0';
                when 3215 => sda_i <= '0';
                when 3216 => sda_i <= '0';
                when 3217 => sda_i <= '0';
                when 3218 => sda_i <= '0';
                when 3219 => sda_i <= '0';
                when 3220 => sda_i <= '0';
                when 3221 => sda_i <= '0';
                when 3222 => sda_i <= '0';
                when 3223 => sda_i <= '0';
                when 3224 => sda_i <= '0';
                when 3225 => sda_i <= '0';
                when 3226 => sda_i <= '0';
                when 3227 => sda_i <= '0';
                when 3228 => sda_i <= '0';
                when 3229 => sda_i <= '0';
                when 3230 => sda_i <= '0';
                when 3231 => sda_i <= '0';
                when 3232 => sda_i <= '0';
                when 3233 => sda_i <= '0';
                when 3234 => sda_i <= '0';
                when 3235 => sda_i <= '0';
                when 3236 => sda_i <= '0';
                when 3237 => sda_i <= '0';
                when 3238 => sda_i <= '1';
                when 3239 => sda_i <= '1';
                when 3240 => sda_i <= '0';
                when 3241 => sda_i <= '0';
                when 3242 => sda_i <= '0';
                when 3243 => sda_i <= '0';
                when 3244 => sda_i <= '0';
                when 3245 => sda_i <= '0';
                when 3246 => sda_i <= '0';
                when 3247 => sda_i <= '0';
                when 3248 => sda_i <= '0';
                when 3249 => sda_i <= '0';
                when 3250 => sda_i <= '0';
                when 3251 => sda_i <= '0';
                when 3252 => sda_i <= '0';
                when 3253 => sda_i <= '0';
                when 3254 => sda_i <= '0';
                when 3255 => sda_i <= '0';
                when 3256 => sda_i <= '0';
                when 3257 => sda_i <= '0';
                when 3258 => sda_i <= '0';
                when 3259 => sda_i <= '0';
                when 3260 => sda_i <= '0';
                when 3261 => sda_i <= '0';
                when 3262 => sda_i <= '0';
                when 3263 => sda_i <= '0';
                when 3264 => sda_i <= '0';
                when 3265 => sda_i <= '0';
                when 3266 => sda_i <= '0';
                when 3267 => sda_i <= '0';
                when 3268 => sda_i <= '0';
                when 3269 => sda_i <= '0';
                when 3270 => sda_i <= '0';
                when 3271 => sda_i <= '0';
                when 3272 => sda_i <= '0';
                when 3273 => sda_i <= '0';
                when 3274 => sda_i <= '0';
                when 3275 => sda_i <= '0';
                when 3276 => sda_i <= '0';
                when 3277 => sda_i <= '0';
                when 3278 => sda_i <= '0';
                when 3279 => sda_i <= '0';
                when 3280 => sda_i <= '0';
                when 3281 => sda_i <= '0';
                when 3282 => sda_i <= '0';
                when 3283 => sda_i <= '0';
                when 3284 => sda_i <= '0';
                when 3285 => sda_i <= '0';
                when 3286 => sda_i <= '0';
                when 3287 => sda_i <= '0';
                when 3288 => sda_i <= '0';
                when 3289 => sda_i <= '0';
                when 3290 => sda_i <= '0';
                when 3291 => sda_i <= '0';
                when 3292 => sda_i <= '0';
                when 3293 => sda_i <= '0';
                when 3294 => sda_i <= '0';
                when 3295 => sda_i <= '0';
                when 3296 => sda_i <= '0';
                when 3297 => sda_i <= '0';
                when 3298 => sda_i <= '0';
                when 3299 => sda_i <= '0';
                when 3300 => sda_i <= '0';
                when 3301 => sda_i <= '0';
                when 3302 => sda_i <= '0';
                when 3303 => sda_i <= '0';
                when 3304 => sda_i <= '0';
                when 3305 => sda_i <= '0';
                when 3306 => sda_i <= '0';
                when 3307 => sda_i <= '0';
                when 3308 => sda_i <= '0';
                when 3309 => sda_i <= '0';
                when 3310 => sda_i <= '0';
                when 3311 => sda_i <= '0';
                when 3312 => sda_i <= '0';
                when 3313 => sda_i <= '0';
                when 3314 => sda_i <= '0';
                when 3315 => sda_i <= '0';
                when 3316 => sda_i <= '0';
                when 3317 => sda_i <= '0';
                when 3318 => sda_i <= '0';
                when 3319 => sda_i <= '0';
                when 3320 => sda_i <= '0';
                when 3321 => sda_i <= '0';
                when 3322 => sda_i <= '0';
                when 3323 => sda_i <= '0';
                when 3324 => sda_i <= '0';
                when 3325 => sda_i <= '0';
                when 3326 => sda_i <= '0';
                when 3327 => sda_i <= '0';
                when 3328 => sda_i <= '0';
                when 3329 => sda_i <= '0';
                when 3330 => sda_i <= '0';
                when 3331 => sda_i <= '0';
                when 3332 => sda_i <= '0';
                when 3333 => sda_i <= '0';
                when 3334 => sda_i <= '0';
                when 3335 => sda_i <= '0';
                when 3336 => sda_i <= '0';
                when 3337 => sda_i <= '0';
                when 3338 => sda_i <= '0';
                when 3339 => sda_i <= '0';
                when 3340 => sda_i <= '0';
                when 3341 => sda_i <= '0';
                when 3342 => sda_i <= '0';
                when 3343 => sda_i <= '0';
                when 3344 => sda_i <= '0';
                when 3345 => sda_i <= '0';
                when 3346 => sda_i <= '1';
                when 3347 => sda_i <= '1';
                when 3348 => sda_i <= '0';
                when 3349 => sda_i <= '0';
                when 3350 => sda_i <= '0';
                when 3351 => sda_i <= '0';
                when 3352 => sda_i <= '0';
                when 3353 => sda_i <= '0';
                when 3354 => sda_i <= '0';
                when 3355 => sda_i <= '0';
                when 3356 => sda_i <= '0';
                when 3357 => sda_i <= '0';
                when 3358 => sda_i <= '0';
                when 3359 => sda_i <= '0';
                when 3360 => sda_i <= '0';
                when 3361 => sda_i <= '0';
                when 3362 => sda_i <= '0';
                when 3363 => sda_i <= '0';
                when 3364 => sda_i <= '0';
                when 3365 => sda_i <= '0';
                when 3366 => sda_i <= '0';
                when 3367 => sda_i <= '0';
                when 3368 => sda_i <= '0';
                when 3369 => sda_i <= '0';
                when 3370 => sda_i <= '0';
                when 3371 => sda_i <= '0';
                when 3372 => sda_i <= '0';
                when 3373 => sda_i <= '0';
                when 3374 => sda_i <= '0';
                when 3375 => sda_i <= '0';
                when 3376 => sda_i <= '0';
                when 3377 => sda_i <= '0';
                when 3378 => sda_i <= '0';
                when 3379 => sda_i <= '0';
                when 3380 => sda_i <= '0';
                when 3381 => sda_i <= '0';
                when 3382 => sda_i <= '0';
                when 3383 => sda_i <= '0';
                when 3384 => sda_i <= '0';
                when 3385 => sda_i <= '0';
                when 3386 => sda_i <= '0';
                when 3387 => sda_i <= '0';
                when 3388 => sda_i <= '0';
                when 3389 => sda_i <= '0';
                when 3390 => sda_i <= '0';
                when 3391 => sda_i <= '0';
                when 3392 => sda_i <= '0';
                when 3393 => sda_i <= '0';
                when 3394 => sda_i <= '0';
                when 3395 => sda_i <= '0';
                when 3396 => sda_i <= '0';
                when 3397 => sda_i <= '0';
                when 3398 => sda_i <= '0';
                when 3399 => sda_i <= '0';
                when 3400 => sda_i <= '0';
                when 3401 => sda_i <= '0';
                when 3402 => sda_i <= '0';
                when 3403 => sda_i <= '0';
                when 3404 => sda_i <= '0';
                when 3405 => sda_i <= '0';
                when 3406 => sda_i <= '0';
                when 3407 => sda_i <= '0';
                when 3408 => sda_i <= '0';
                when 3409 => sda_i <= '0';
                when 3410 => sda_i <= '0';
                when 3411 => sda_i <= '0';
                when 3412 => sda_i <= '0';
                when 3413 => sda_i <= '0';
                when 3414 => sda_i <= '0';
                when 3415 => sda_i <= '0';
                when 3416 => sda_i <= '0';
                when 3417 => sda_i <= '0';
                when 3418 => sda_i <= '0';
                when 3419 => sda_i <= '0';
                when 3420 => sda_i <= '0';
                when 3421 => sda_i <= '0';
                when 3422 => sda_i <= '0';
                when 3423 => sda_i <= '0';
                when 3424 => sda_i <= '0';
                when 3425 => sda_i <= '0';
                when 3426 => sda_i <= '0';
                when 3427 => sda_i <= '0';
                when 3428 => sda_i <= '0';
                when 3429 => sda_i <= '0';
                when 3430 => sda_i <= '0';
                when 3431 => sda_i <= '0';
                when 3432 => sda_i <= '0';
                when 3433 => sda_i <= '0';
                when 3434 => sda_i <= '0';
                when 3435 => sda_i <= '0';
                when 3436 => sda_i <= '0';
                when 3437 => sda_i <= '0';
                when 3438 => sda_i <= '0';
                when 3439 => sda_i <= '0';
                when 3440 => sda_i <= '0';
                when 3441 => sda_i <= '0';
                when 3442 => sda_i <= '0';
                when 3443 => sda_i <= '0';
                when 3444 => sda_i <= '0';
                when 3445 => sda_i <= '0';
                when 3446 => sda_i <= '0';
                when 3447 => sda_i <= '0';
                when 3448 => sda_i <= '0';
                when 3449 => sda_i <= '0';
                when 3450 => sda_i <= '0';
                when 3451 => sda_i <= '0';
                when 3452 => sda_i <= '0';
                when 3453 => sda_i <= '0';
                when 3454 => sda_i <= '1';
                when 3455 => sda_i <= '1';
                when 3456 => sda_i <= '0';
                when 3457 => sda_i <= '0';
                when 3458 => sda_i <= '0';
                when 3459 => sda_i <= '0';
                when 3460 => sda_i <= '0';
                when 3461 => sda_i <= '0';
                when 3462 => sda_i <= '0';
                when 3463 => sda_i <= '0';
                when 3464 => sda_i <= '0';
                when 3465 => sda_i <= '0';
                when 3466 => sda_i <= '0';
                when 3467 => sda_i <= '0';
                when 3468 => sda_i <= '0';
                when 3469 => sda_i <= '0';
                when 3470 => sda_i <= '0';
                when 3471 => sda_i <= '0';
                when 3472 => sda_i <= '0';
                when 3473 => sda_i <= '0';
                when 3474 => sda_i <= '0';
                when 3475 => sda_i <= '0';
                when 3476 => sda_i <= '0';
                when 3477 => sda_i <= '0';
                when 3478 => sda_i <= '0';
                when 3479 => sda_i <= '0';
                when 3480 => sda_i <= '0';
                when 3481 => sda_i <= '0';
                when 3482 => sda_i <= '0';
                when 3483 => sda_i <= '0';
                when 3484 => sda_i <= '0';
                when 3485 => sda_i <= '0';
                when 3486 => sda_i <= '0';
                when 3487 => sda_i <= '0';
                when 3488 => sda_i <= '0';
                when 3489 => sda_i <= '0';
                when 3490 => sda_i <= '0';
                when 3491 => sda_i <= '0';
                when 3492 => sda_i <= '0';
                when 3493 => sda_i <= '0';
                when 3494 => sda_i <= '0';
                when 3495 => sda_i <= '0';
                when 3496 => sda_i <= '0';
                when 3497 => sda_i <= '0';
                when 3498 => sda_i <= '0';
                when 3499 => sda_i <= '0';
                when 3500 => sda_i <= '0';
                when 3501 => sda_i <= '0';
                when 3502 => sda_i <= '0';
                when 3503 => sda_i <= '0';
                when 3504 => sda_i <= '0';
                when 3505 => sda_i <= '0';
                when 3506 => sda_i <= '0';
                when 3507 => sda_i <= '0';
                when 3508 => sda_i <= '0';
                when 3509 => sda_i <= '0';
                when 3510 => sda_i <= '0';
                when 3511 => sda_i <= '0';
                when 3512 => sda_i <= '0';
                when 3513 => sda_i <= '0';
                when 3514 => sda_i <= '0';
                when 3515 => sda_i <= '0';
                when 3516 => sda_i <= '0';
                when 3517 => sda_i <= '0';
                when 3518 => sda_i <= '0';
                when 3519 => sda_i <= '0';
                when 3520 => sda_i <= '0';
                when 3521 => sda_i <= '0';
                when 3522 => sda_i <= '0';
                when 3523 => sda_i <= '0';
                when 3524 => sda_i <= '0';
                when 3525 => sda_i <= '0';
                when 3526 => sda_i <= '0';
                when 3527 => sda_i <= '0';
                when 3528 => sda_i <= '0';
                when 3529 => sda_i <= '0';
                when 3530 => sda_i <= '0';
                when 3531 => sda_i <= '0';
                when 3532 => sda_i <= '0';
                when 3533 => sda_i <= '0';
                when 3534 => sda_i <= '0';
                when 3535 => sda_i <= '0';
                when 3536 => sda_i <= '0';
                when 3537 => sda_i <= '0';
                when 3538 => sda_i <= '0';
                when 3539 => sda_i <= '0';
                when 3540 => sda_i <= '0';
                when 3541 => sda_i <= '0';
                when 3542 => sda_i <= '0';
                when 3543 => sda_i <= '0';
                when 3544 => sda_i <= '0';
                when 3545 => sda_i <= '0';
                when 3546 => sda_i <= '0';
                when 3547 => sda_i <= '0';
                when 3548 => sda_i <= '0';
                when 3549 => sda_i <= '0';
                when 3550 => sda_i <= '0';
                when 3551 => sda_i <= '0';
                when 3552 => sda_i <= '0';
                when 3553 => sda_i <= '0';
                when 3554 => sda_i <= '0';
                when 3555 => sda_i <= '0';
                when 3556 => sda_i <= '0';
                when 3557 => sda_i <= '0';
                when 3558 => sda_i <= '0';
                when 3559 => sda_i <= '0';
                when 3560 => sda_i <= '0';
                when 3561 => sda_i <= '0';
                when 3562 => sda_i <= '1';
                when 3563 => sda_i <= '1';
                when 3564 => sda_i <= '0';
                when 3565 => sda_i <= '0';
                when 3566 => sda_i <= '0';
                when 3567 => sda_i <= '0';
                when 3568 => sda_i <= '0';
                when 3569 => sda_i <= '0';
                when 3570 => sda_i <= '0';
                when 3571 => sda_i <= '0';
                when 3572 => sda_i <= '0';
                when 3573 => sda_i <= '0';
                when 3574 => sda_i <= '0';
                when 3575 => sda_i <= '0';
                when 3576 => sda_i <= '0';
                when 3577 => sda_i <= '0';
                when 3578 => sda_i <= '0';
                when 3579 => sda_i <= '0';
                when 3580 => sda_i <= '0';
                when 3581 => sda_i <= '0';
                when 3582 => sda_i <= '0';
                when 3583 => sda_i <= '0';
                when 3584 => sda_i <= '0';
                when 3585 => sda_i <= '0';
                when 3586 => sda_i <= '0';
                when 3587 => sda_i <= '0';
                when 3588 => sda_i <= '0';
                when 3589 => sda_i <= '0';
                when 3590 => sda_i <= '0';
                when 3591 => sda_i <= '0';
                when 3592 => sda_i <= '0';
                when 3593 => sda_i <= '0';
                when 3594 => sda_i <= '0';
                when 3595 => sda_i <= '0';
                when 3596 => sda_i <= '0';
                when 3597 => sda_i <= '0';
                when 3598 => sda_i <= '0';
                when 3599 => sda_i <= '0';
                when 3600 => sda_i <= '0';
                when 3601 => sda_i <= '0';
                when 3602 => sda_i <= '0';
                when 3603 => sda_i <= '0';
                when 3604 => sda_i <= '0';
                when 3605 => sda_i <= '0';
                when 3606 => sda_i <= '0';
                when 3607 => sda_i <= '0';
                when 3608 => sda_i <= '0';
                when 3609 => sda_i <= '0';
                when 3610 => sda_i <= '0';
                when 3611 => sda_i <= '0';
                when 3612 => sda_i <= '0';
                when 3613 => sda_i <= '0';
                when 3614 => sda_i <= '0';
                when 3615 => sda_i <= '0';
                when 3616 => sda_i <= '0';
                when 3617 => sda_i <= '0';
                when 3618 => sda_i <= '0';
                when 3619 => sda_i <= '0';
                when 3620 => sda_i <= '0';
                when 3621 => sda_i <= '0';
                when 3622 => sda_i <= '0';
                when 3623 => sda_i <= '0';
                when 3624 => sda_i <= '0';
                when 3625 => sda_i <= '0';
                when 3626 => sda_i <= '0';
                when 3627 => sda_i <= '0';
                when 3628 => sda_i <= '0';
                when 3629 => sda_i <= '0';
                when 3630 => sda_i <= '0';
                when 3631 => sda_i <= '0';
                when 3632 => sda_i <= '0';
                when 3633 => sda_i <= '0';
                when 3634 => sda_i <= '0';
                when 3635 => sda_i <= '0';
                when 3636 => sda_i <= '0';
                when 3637 => sda_i <= '0';
                when 3638 => sda_i <= '0';
                when 3639 => sda_i <= '0';
                when 3640 => sda_i <= '0';
                when 3641 => sda_i <= '0';
                when 3642 => sda_i <= '0';
                when 3643 => sda_i <= '0';
                when 3644 => sda_i <= '0';
                when 3645 => sda_i <= '0';
                when 3646 => sda_i <= '0';
                when 3647 => sda_i <= '0';
                when 3648 => sda_i <= '0';
                when 3649 => sda_i <= '0';
                when 3650 => sda_i <= '0';
                when 3651 => sda_i <= '0';
                when 3652 => sda_i <= '0';
                when 3653 => sda_i <= '0';
                when 3654 => sda_i <= '0';
                when 3655 => sda_i <= '0';
                when 3656 => sda_i <= '0';
                when 3657 => sda_i <= '0';
                when 3658 => sda_i <= '0';
                when 3659 => sda_i <= '0';
                when 3660 => sda_i <= '0';
                when 3661 => sda_i <= '0';
                when 3662 => sda_i <= '0';
                when 3663 => sda_i <= '0';
                when 3664 => sda_i <= '0';
                when 3665 => sda_i <= '0';
                when 3666 => sda_i <= '0';
                when 3667 => sda_i <= '0';
                when 3668 => sda_i <= '0';
                when 3669 => sda_i <= '0';
                when 3670 => sda_i <= '1';
                when 3671 => sda_i <= '1';
                when 3672 => sda_i <= '0';
                when 3673 => sda_i <= '0';
                when 3674 => sda_i <= '0';
                when 3675 => sda_i <= '0';
                when 3676 => sda_i <= '0';
                when 3677 => sda_i <= '0';
                when 3678 => sda_i <= '0';
                when 3679 => sda_i <= '0';
                when 3680 => sda_i <= '0';
                when 3681 => sda_i <= '0';
                when 3682 => sda_i <= '0';
                when 3683 => sda_i <= '0';
                when 3684 => sda_i <= '0';
                when 3685 => sda_i <= '0';
                when 3686 => sda_i <= '0';
                when 3687 => sda_i <= '0';
                when 3688 => sda_i <= '0';
                when 3689 => sda_i <= '0';
                when 3690 => sda_i <= '0';
                when 3691 => sda_i <= '0';
                when 3692 => sda_i <= '0';
                when 3693 => sda_i <= '0';
                when 3694 => sda_i <= '0';
                when 3695 => sda_i <= '0';
                when 3696 => sda_i <= '0';
                when 3697 => sda_i <= '0';
                when 3698 => sda_i <= '0';
                when 3699 => sda_i <= '0';
                when 3700 => sda_i <= '0';
                when 3701 => sda_i <= '0';
                when 3702 => sda_i <= '0';
                when 3703 => sda_i <= '0';
                when 3704 => sda_i <= '0';
                when 3705 => sda_i <= '0';
                when 3706 => sda_i <= '0';
                when 3707 => sda_i <= '0';
                when 3708 => sda_i <= '0';
                when 3709 => sda_i <= '0';
                when 3710 => sda_i <= '0';
                when 3711 => sda_i <= '0';
                when 3712 => sda_i <= '0';
                when 3713 => sda_i <= '0';
                when 3714 => sda_i <= '0';
                when 3715 => sda_i <= '0';
                when 3716 => sda_i <= '0';
                when 3717 => sda_i <= '0';
                when 3718 => sda_i <= '0';
                when 3719 => sda_i <= '0';
                when 3720 => sda_i <= '0';
                when 3721 => sda_i <= '0';
                when 3722 => sda_i <= '0';
                when 3723 => sda_i <= '0';
                when 3724 => sda_i <= '0';
                when 3725 => sda_i <= '0';
                when 3726 => sda_i <= '0';
                when 3727 => sda_i <= '0';
                when 3728 => sda_i <= '0';
                when 3729 => sda_i <= '0';
                when 3730 => sda_i <= '0';
                when 3731 => sda_i <= '0';
                when 3732 => sda_i <= '0';
                when 3733 => sda_i <= '0';
                when 3734 => sda_i <= '0';
                when 3735 => sda_i <= '0';
                when 3736 => sda_i <= '0';
                when 3737 => sda_i <= '0';
                when 3738 => sda_i <= '0';
                when 3739 => sda_i <= '0';
                when 3740 => sda_i <= '0';
                when 3741 => sda_i <= '0';
                when 3742 => sda_i <= '0';
                when 3743 => sda_i <= '0';
                when 3744 => sda_i <= '0';
                when 3745 => sda_i <= '0';
                when 3746 => sda_i <= '0';
                when 3747 => sda_i <= '0';
                when 3748 => sda_i <= '0';
                when 3749 => sda_i <= '0';
                when 3750 => sda_i <= '0';
                when 3751 => sda_i <= '0';
                when 3752 => sda_i <= '0';
                when 3753 => sda_i <= '0';
                when 3754 => sda_i <= '0';
                when 3755 => sda_i <= '0';
                when 3756 => sda_i <= '0';
                when 3757 => sda_i <= '0';
                when 3758 => sda_i <= '0';
                when 3759 => sda_i <= '0';
                when 3760 => sda_i <= '0';
                when 3761 => sda_i <= '0';
                when 3762 => sda_i <= '0';
                when 3763 => sda_i <= '0';
                when 3764 => sda_i <= '0';
                when 3765 => sda_i <= '0';
                when 3766 => sda_i <= '0';
                when 3767 => sda_i <= '0';
                when 3768 => sda_i <= '0';
                when 3769 => sda_i <= '0';
                when 3770 => sda_i <= '0';
                when 3771 => sda_i <= '0';
                when 3772 => sda_i <= '0';
                when 3773 => sda_i <= '0';
                when 3774 => sda_i <= '0';
                when 3775 => sda_i <= '0';
                when 3776 => sda_i <= '0';
                when 3777 => sda_i <= '0';
                when 3778 => sda_i <= '1';
                when 3779 => sda_i <= '1';
                when 3780 => sda_i <= '0';
                when 3781 => sda_i <= '0';
                when 3782 => sda_i <= '0';
                when 3783 => sda_i <= '0';
                when 3784 => sda_i <= '0';
                when 3785 => sda_i <= '0';
                when 3786 => sda_i <= '0';
                when 3787 => sda_i <= '0';
                when 3788 => sda_i <= '0';
                when 3789 => sda_i <= '0';
                when 3790 => sda_i <= '0';
                when 3791 => sda_i <= '0';
                when 3792 => sda_i <= '0';
                when 3793 => sda_i <= '0';
                when 3794 => sda_i <= '0';
                when 3795 => sda_i <= '0';
                when 3796 => sda_i <= '0';
                when 3797 => sda_i <= '0';
                when 3798 => sda_i <= '0';
                when 3799 => sda_i <= '0';
                when 3800 => sda_i <= '0';
                when 3801 => sda_i <= '0';
                when 3802 => sda_i <= '0';
                when 3803 => sda_i <= '0';
                when 3804 => sda_i <= '0';
                when 3805 => sda_i <= '0';
                when 3806 => sda_i <= '0';
                when 3807 => sda_i <= '0';
                when 3808 => sda_i <= '0';
                when 3809 => sda_i <= '0';
                when 3810 => sda_i <= '0';
                when 3811 => sda_i <= '0';
                when 3812 => sda_i <= '0';
                when 3813 => sda_i <= '0';
                when 3814 => sda_i <= '0';
                when 3815 => sda_i <= '0';
                when 3816 => sda_i <= '0';
                when 3817 => sda_i <= '0';
                when 3818 => sda_i <= '0';
                when 3819 => sda_i <= '0';
                when 3820 => sda_i <= '0';
                when 3821 => sda_i <= '0';
                when 3822 => sda_i <= '0';
                when 3823 => sda_i <= '0';
                when 3824 => sda_i <= '0';
                when 3825 => sda_i <= '0';
                when 3826 => sda_i <= '0';
                when 3827 => sda_i <= '0';
                when 3828 => sda_i <= '0';
                when 3829 => sda_i <= '0';
                when 3830 => sda_i <= '0';
                when 3831 => sda_i <= '0';
                when 3832 => sda_i <= '0';
                when 3833 => sda_i <= '0';
                when 3834 => sda_i <= '0';
                when 3835 => sda_i <= '0';
                when 3836 => sda_i <= '0';
                when 3837 => sda_i <= '0';
                when 3838 => sda_i <= '0';
                when 3839 => sda_i <= '0';
                when 3840 => sda_i <= '0';
                when 3841 => sda_i <= '0';
                when 3842 => sda_i <= '0';
                when 3843 => sda_i <= '0';
                when 3844 => sda_i <= '0';
                when 3845 => sda_i <= '0';
                when 3846 => sda_i <= '0';
                when 3847 => sda_i <= '0';
                when 3848 => sda_i <= '0';
                when 3849 => sda_i <= '0';
                when 3850 => sda_i <= '0';
                when 3851 => sda_i <= '0';
                when 3852 => sda_i <= '0';
                when 3853 => sda_i <= '0';
                when 3854 => sda_i <= '0';
                when 3855 => sda_i <= '0';
                when 3856 => sda_i <= '0';
                when 3857 => sda_i <= '0';
                when 3858 => sda_i <= '0';
                when 3859 => sda_i <= '0';
                when 3860 => sda_i <= '0';
                when 3861 => sda_i <= '0';
                when 3862 => sda_i <= '0';
                when 3863 => sda_i <= '0';
                when 3864 => sda_i <= '0';
                when 3865 => sda_i <= '0';
                when 3866 => sda_i <= '0';
                when 3867 => sda_i <= '0';
                when 3868 => sda_i <= '0';
                when 3869 => sda_i <= '0';
                when 3870 => sda_i <= '0';
                when 3871 => sda_i <= '0';
                when 3872 => sda_i <= '0';
                when 3873 => sda_i <= '0';
                when 3874 => sda_i <= '0';
                when 3875 => sda_i <= '0';
                when 3876 => sda_i <= '0';
                when 3877 => sda_i <= '0';
                when 3878 => sda_i <= '0';
                when 3879 => sda_i <= '0';
                when 3880 => sda_i <= '0';
                when 3881 => sda_i <= '0';
                when 3882 => sda_i <= '0';
                when 3883 => sda_i <= '0';
                when 3884 => sda_i <= '0';
                when 3885 => sda_i <= '0';
                when 3886 => sda_i <= '1';
                when 3887 => sda_i <= '1';
                when 3888 => sda_i <= '0';
                when 3889 => sda_i <= '0';
                when 3890 => sda_i <= '0';
                when 3891 => sda_i <= '0';
                when 3892 => sda_i <= '0';
                when 3893 => sda_i <= '0';
                when 3894 => sda_i <= '0';
                when 3895 => sda_i <= '0';
                when 3896 => sda_i <= '0';
                when 3897 => sda_i <= '0';
                when 3898 => sda_i <= '0';
                when 3899 => sda_i <= '0';
                when 3900 => sda_i <= '0';
                when 3901 => sda_i <= '0';
                when 3902 => sda_i <= '0';
                when 3903 => sda_i <= '0';
                when 3904 => sda_i <= '0';
                when 3905 => sda_i <= '0';
                when 3906 => sda_i <= '0';
                when 3907 => sda_i <= '0';
                when 3908 => sda_i <= '0';
                when 3909 => sda_i <= '0';
                when 3910 => sda_i <= '0';
                when 3911 => sda_i <= '0';
                when 3912 => sda_i <= '0';
                when 3913 => sda_i <= '0';
                when 3914 => sda_i <= '0';
                when 3915 => sda_i <= '0';
                when 3916 => sda_i <= '0';
                when 3917 => sda_i <= '0';
                when 3918 => sda_i <= '0';
                when 3919 => sda_i <= '0';
                when 3920 => sda_i <= '0';
                when 3921 => sda_i <= '0';
                when 3922 => sda_i <= '0';
                when 3923 => sda_i <= '0';
                when 3924 => sda_i <= '0';
                when 3925 => sda_i <= '0';
                when 3926 => sda_i <= '0';
                when 3927 => sda_i <= '0';
                when 3928 => sda_i <= '0';
                when 3929 => sda_i <= '0';
                when 3930 => sda_i <= '0';
                when 3931 => sda_i <= '0';
                when 3932 => sda_i <= '0';
                when 3933 => sda_i <= '0';
                when 3934 => sda_i <= '0';
                when 3935 => sda_i <= '0';
                when 3936 => sda_i <= '0';
                when 3937 => sda_i <= '0';
                when 3938 => sda_i <= '0';
                when 3939 => sda_i <= '0';
                when 3940 => sda_i <= '0';
                when 3941 => sda_i <= '0';
                when 3942 => sda_i <= '0';
                when 3943 => sda_i <= '0';
                when 3944 => sda_i <= '0';
                when 3945 => sda_i <= '0';
                when 3946 => sda_i <= '0';
                when 3947 => sda_i <= '0';
                when 3948 => sda_i <= '0';
                when 3949 => sda_i <= '0';
                when 3950 => sda_i <= '0';
                when 3951 => sda_i <= '0';
                when 3952 => sda_i <= '0';
                when 3953 => sda_i <= '0';
                when 3954 => sda_i <= '0';
                when 3955 => sda_i <= '0';
                when 3956 => sda_i <= '0';
                when 3957 => sda_i <= '0';
                when 3958 => sda_i <= '0';
                when 3959 => sda_i <= '0';
                when 3960 => sda_i <= '0';
                when 3961 => sda_i <= '0';
                when 3962 => sda_i <= '0';
                when 3963 => sda_i <= '0';
                when 3964 => sda_i <= '0';
                when 3965 => sda_i <= '0';
                when 3966 => sda_i <= '0';
                when 3967 => sda_i <= '0';
                when 3968 => sda_i <= '0';
                when 3969 => sda_i <= '0';
                when 3970 => sda_i <= '0';
                when 3971 => sda_i <= '0';
                when 3972 => sda_i <= '0';
                when 3973 => sda_i <= '0';
                when 3974 => sda_i <= '0';
                when 3975 => sda_i <= '0';
                when 3976 => sda_i <= '0';
                when 3977 => sda_i <= '0';
                when 3978 => sda_i <= '0';
                when 3979 => sda_i <= '0';
                when 3980 => sda_i <= '0';
                when 3981 => sda_i <= '0';
                when 3982 => sda_i <= '0';
                when 3983 => sda_i <= '0';
                when 3984 => sda_i <= '0';
                when 3985 => sda_i <= '0';
                when 3986 => sda_i <= '0';
                when 3987 => sda_i <= '0';
                when 3988 => sda_i <= '0';
                when 3989 => sda_i <= '0';
                when 3990 => sda_i <= '0';
                when 3991 => sda_i <= '0';
                when 3992 => sda_i <= '0';
                when 3993 => sda_i <= '0';
                when 3994 => sda_i <= '1';
                when 3995 => sda_i <= '1';
                when 3996 => sda_i <= '0';
                when 3997 => sda_i <= '0';
                when 3998 => sda_i <= '0';
                when 3999 => sda_i <= '0';
                when 4000 => sda_i <= '0';
                when 4001 => sda_i <= '0';
                when 4002 => sda_i <= '0';
                when 4003 => sda_i <= '0';
                when 4004 => sda_i <= '0';
                when 4005 => sda_i <= '0';
                when 4006 => sda_i <= '0';
                when 4007 => sda_i <= '0';
                when 4008 => sda_i <= '0';
                when 4009 => sda_i <= '0';
                when 4010 => sda_i <= '0';
                when 4011 => sda_i <= '0';
                when 4012 => sda_i <= '0';
                when 4013 => sda_i <= '0';
                when 4014 => sda_i <= '0';
                when 4015 => sda_i <= '0';
                when 4016 => sda_i <= '0';
                when 4017 => sda_i <= '0';
                when 4018 => sda_i <= '0';
                when 4019 => sda_i <= '0';
                when 4020 => sda_i <= '0';
                when 4021 => sda_i <= '0';
                when 4022 => sda_i <= '0';
                when 4023 => sda_i <= '0';
                when 4024 => sda_i <= '0';
                when 4025 => sda_i <= '0';
                when 4026 => sda_i <= '0';
                when 4027 => sda_i <= '0';
                when 4028 => sda_i <= '0';
                when 4029 => sda_i <= '0';
                when 4030 => sda_i <= '0';
                when 4031 => sda_i <= '0';
                when 4032 => sda_i <= '0';
                when 4033 => sda_i <= '0';
                when 4034 => sda_i <= '0';
                when 4035 => sda_i <= '0';
                when 4036 => sda_i <= '0';
                when 4037 => sda_i <= '0';
                when 4038 => sda_i <= '0';
                when 4039 => sda_i <= '0';
                when 4040 => sda_i <= '0';
                when 4041 => sda_i <= '0';
                when 4042 => sda_i <= '0';
                when 4043 => sda_i <= '0';
                when 4044 => sda_i <= '0';
                when 4045 => sda_i <= '0';
                when 4046 => sda_i <= '0';
                when 4047 => sda_i <= '0';
                when 4048 => sda_i <= '0';
                when 4049 => sda_i <= '0';
                when 4050 => sda_i <= '0';
                when 4051 => sda_i <= '0';
                when 4052 => sda_i <= '0';
                when 4053 => sda_i <= '0';
                when 4054 => sda_i <= '0';
                when 4055 => sda_i <= '0';
                when 4056 => sda_i <= '0';
                when 4057 => sda_i <= '0';
                when 4058 => sda_i <= '0';
                when 4059 => sda_i <= '0';
                when 4060 => sda_i <= '0';
                when 4061 => sda_i <= '0';
                when 4062 => sda_i <= '0';
                when 4063 => sda_i <= '0';
                when 4064 => sda_i <= '0';
                when 4065 => sda_i <= '0';
                when 4066 => sda_i <= '0';
                when 4067 => sda_i <= '0';
                when 4068 => sda_i <= '0';
                when 4069 => sda_i <= '0';
                when 4070 => sda_i <= '0';
                when 4071 => sda_i <= '0';
                when 4072 => sda_i <= '0';
                when 4073 => sda_i <= '0';
                when 4074 => sda_i <= '0';
                when 4075 => sda_i <= '0';
                when 4076 => sda_i <= '0';
                when 4077 => sda_i <= '0';
                when 4078 => sda_i <= '0';
                when 4079 => sda_i <= '0';
                when 4080 => sda_i <= '0';
                when 4081 => sda_i <= '0';
                when 4082 => sda_i <= '0';
                when 4083 => sda_i <= '0';
                when 4084 => sda_i <= '0';
                when 4085 => sda_i <= '0';
                when 4086 => sda_i <= '0';
                when 4087 => sda_i <= '0';
                when 4088 => sda_i <= '0';
                when 4089 => sda_i <= '0';
                when 4090 => sda_i <= '0';
                when 4091 => sda_i <= '0';
                when 4092 => sda_i <= '0';
                when 4093 => sda_i <= '0';
                when 4094 => sda_i <= '0';
                when 4095 => sda_i <= '0';
                when 4096 => sda_i <= '0';
                when 4097 => sda_i <= '0';
                when 4098 => sda_i <= '0';
                when 4099 => sda_i <= '0';
                when 4100 => sda_i <= '0';
                when 4101 => sda_i <= '0';
                when 4102 => sda_i <= '1';
                when 4103 => sda_i <= '1';
                when 4104 => sda_i <= '0';
                when 4105 => sda_i <= '0';
                when 4106 => sda_i <= '0';
                when 4107 => sda_i <= '0';
                when 4108 => sda_i <= '0';
                when 4109 => sda_i <= '0';
                when 4110 => sda_i <= '0';
                when 4111 => sda_i <= '0';
                when 4112 => sda_i <= '0';
                when 4113 => sda_i <= '0';
                when 4114 => sda_i <= '0';
                when 4115 => sda_i <= '0';
                when 4116 => sda_i <= '0';
                when 4117 => sda_i <= '0';
                when 4118 => sda_i <= '0';
                when 4119 => sda_i <= '0';
                when 4120 => sda_i <= '0';
                when 4121 => sda_i <= '0';
                when 4122 => sda_i <= '0';
                when 4123 => sda_i <= '0';
                when 4124 => sda_i <= '0';
                when 4125 => sda_i <= '0';
                when 4126 => sda_i <= '0';
                when 4127 => sda_i <= '0';
                when 4128 => sda_i <= '0';
                when 4129 => sda_i <= '0';
                when 4130 => sda_i <= '0';
                when 4131 => sda_i <= '0';
                when 4132 => sda_i <= '0';
                when 4133 => sda_i <= '0';
                when 4134 => sda_i <= '0';
                when 4135 => sda_i <= '0';
                when 4136 => sda_i <= '0';
                when 4137 => sda_i <= '0';
                when 4138 => sda_i <= '0';
                when 4139 => sda_i <= '0';
                when 4140 => sda_i <= '0';
                when 4141 => sda_i <= '0';
                when 4142 => sda_i <= '0';
                when 4143 => sda_i <= '0';
                when 4144 => sda_i <= '0';
                when 4145 => sda_i <= '0';
                when 4146 => sda_i <= '0';
                when 4147 => sda_i <= '0';
                when 4148 => sda_i <= '0';
                when 4149 => sda_i <= '0';
                when 4150 => sda_i <= '0';
                when 4151 => sda_i <= '0';
                when 4152 => sda_i <= '0';
                when 4153 => sda_i <= '0';
                when 4154 => sda_i <= '0';
                when 4155 => sda_i <= '0';
                when 4156 => sda_i <= '0';
                when 4157 => sda_i <= '0';
                when 4158 => sda_i <= '0';
                when 4159 => sda_i <= '0';
                when 4160 => sda_i <= '0';
                when 4161 => sda_i <= '0';
                when 4162 => sda_i <= '0';
                when 4163 => sda_i <= '0';
                when 4164 => sda_i <= '0';
                when 4165 => sda_i <= '0';
                when 4166 => sda_i <= '0';
                when 4167 => sda_i <= '0';
                when 4168 => sda_i <= '0';
                when 4169 => sda_i <= '0';
                when 4170 => sda_i <= '0';
                when 4171 => sda_i <= '0';
                when 4172 => sda_i <= '0';
                when 4173 => sda_i <= '0';
                when 4174 => sda_i <= '0';
                when 4175 => sda_i <= '0';
                when 4176 => sda_i <= '0';
                when 4177 => sda_i <= '0';
                when 4178 => sda_i <= '0';
                when 4179 => sda_i <= '0';
                when 4180 => sda_i <= '0';
                when 4181 => sda_i <= '0';
                when 4182 => sda_i <= '0';
                when 4183 => sda_i <= '0';
                when 4184 => sda_i <= '0';
                when 4185 => sda_i <= '0';
                when 4186 => sda_i <= '0';
                when 4187 => sda_i <= '0';
                when 4188 => sda_i <= '0';
                when 4189 => sda_i <= '0';
                when 4190 => sda_i <= '0';
                when 4191 => sda_i <= '0';
                when 4192 => sda_i <= '0';
                when 4193 => sda_i <= '0';
                when 4194 => sda_i <= '0';
                when 4195 => sda_i <= '0';
                when 4196 => sda_i <= '0';
                when 4197 => sda_i <= '0';
                when 4198 => sda_i <= '0';
                when 4199 => sda_i <= '0';
                when 4200 => sda_i <= '0';
                when 4201 => sda_i <= '0';
                when 4202 => sda_i <= '0';
                when 4203 => sda_i <= '0';
                when 4204 => sda_i <= '0';
                when 4205 => sda_i <= '0';
                when 4206 => sda_i <= '0';
                when 4207 => sda_i <= '0';
                when 4208 => sda_i <= '0';
                when 4209 => sda_i <= '0';
                when 4210 => sda_i <= '1';
                when 4211 => sda_i <= '1';
                when 4212 => sda_i <= '0';
                when 4213 => sda_i <= '0';
                when 4214 => sda_i <= '0';
                when 4215 => sda_i <= '0';
                when 4216 => sda_i <= '0';
                when 4217 => sda_i <= '0';
                when 4218 => sda_i <= '0';
                when 4219 => sda_i <= '0';
                when 4220 => sda_i <= '0';
                when 4221 => sda_i <= '0';
                when 4222 => sda_i <= '0';
                when 4223 => sda_i <= '0';
                when 4224 => sda_i <= '0';
                when 4225 => sda_i <= '0';
                when 4226 => sda_i <= '0';
                when 4227 => sda_i <= '0';
                when 4228 => sda_i <= '0';
                when 4229 => sda_i <= '0';
                when 4230 => sda_i <= '0';
                when 4231 => sda_i <= '0';
                when 4232 => sda_i <= '0';
                when 4233 => sda_i <= '0';
                when 4234 => sda_i <= '0';
                when 4235 => sda_i <= '0';
                when 4236 => sda_i <= '0';
                when 4237 => sda_i <= '0';
                when 4238 => sda_i <= '0';
                when 4239 => sda_i <= '0';
                when 4240 => sda_i <= '0';
                when 4241 => sda_i <= '0';
                when 4242 => sda_i <= '0';
                when 4243 => sda_i <= '0';
                when 4244 => sda_i <= '0';
                when 4245 => sda_i <= '0';
                when 4246 => sda_i <= '0';
                when 4247 => sda_i <= '0';
                when 4248 => sda_i <= '0';
                when 4249 => sda_i <= '0';
                when 4250 => sda_i <= '0';
                when 4251 => sda_i <= '0';
                when 4252 => sda_i <= '0';
                when 4253 => sda_i <= '0';
                when 4254 => sda_i <= '0';
                when 4255 => sda_i <= '0';
                when 4256 => sda_i <= '0';
                when 4257 => sda_i <= '0';
                when 4258 => sda_i <= '0';
                when 4259 => sda_i <= '0';
                when 4260 => sda_i <= '0';
                when 4261 => sda_i <= '0';
                when 4262 => sda_i <= '0';
                when 4263 => sda_i <= '0';
                when 4264 => sda_i <= '0';
                when 4265 => sda_i <= '0';
                when 4266 => sda_i <= '0';
                when 4267 => sda_i <= '0';
                when 4268 => sda_i <= '0';
                when 4269 => sda_i <= '0';
                when 4270 => sda_i <= '0';
                when 4271 => sda_i <= '0';
                when 4272 => sda_i <= '0';
                when 4273 => sda_i <= '0';
                when 4274 => sda_i <= '0';
                when 4275 => sda_i <= '0';
                when 4276 => sda_i <= '0';
                when 4277 => sda_i <= '0';
                when 4278 => sda_i <= '0';
                when 4279 => sda_i <= '0';
                when 4280 => sda_i <= '0';
                when 4281 => sda_i <= '0';
                when 4282 => sda_i <= '0';
                when 4283 => sda_i <= '0';
                when 4284 => sda_i <= '0';
                when 4285 => sda_i <= '0';
                when 4286 => sda_i <= '0';
                when 4287 => sda_i <= '0';
                when 4288 => sda_i <= '0';
                when 4289 => sda_i <= '0';
                when 4290 => sda_i <= '0';
                when 4291 => sda_i <= '0';
                when 4292 => sda_i <= '0';
                when 4293 => sda_i <= '0';
                when 4294 => sda_i <= '0';
                when 4295 => sda_i <= '0';
                when 4296 => sda_i <= '0';
                when 4297 => sda_i <= '0';
                when 4298 => sda_i <= '0';
                when 4299 => sda_i <= '0';
                when 4300 => sda_i <= '0';
                when 4301 => sda_i <= '0';
                when 4302 => sda_i <= '0';
                when 4303 => sda_i <= '0';
                when 4304 => sda_i <= '0';
                when 4305 => sda_i <= '0';
                when 4306 => sda_i <= '0';
                when 4307 => sda_i <= '0';
                when 4308 => sda_i <= '0';
                when 4309 => sda_i <= '0';
                when 4310 => sda_i <= '0';
                when 4311 => sda_i <= '0';
                when 4312 => sda_i <= '0';
                when 4313 => sda_i <= '0';
                when 4314 => sda_i <= '0';
                when 4315 => sda_i <= '0';
                when 4316 => sda_i <= '0';
                when 4317 => sda_i <= '0';
                when 4318 => sda_i <= '1';
                when 4319 => sda_i <= '1';
                when 4320 => sda_i <= '0';
                when 4321 => sda_i <= '0';
                when 4322 => sda_i <= '0';
                when 4323 => sda_i <= '0';
                when 4324 => sda_i <= '0';
                when 4325 => sda_i <= '0';
                when 4326 => sda_i <= '0';
                when 4327 => sda_i <= '0';
                when 4328 => sda_i <= '0';
                when 4329 => sda_i <= '0';
                when 4330 => sda_i <= '0';
                when 4331 => sda_i <= '0';
                when 4332 => sda_i <= '0';
                when 4333 => sda_i <= '0';
                when 4334 => sda_i <= '0';
                when 4335 => sda_i <= '0';
                when 4336 => sda_i <= '0';
                when 4337 => sda_i <= '0';
                when 4338 => sda_i <= '0';
                when 4339 => sda_i <= '0';
                when 4340 => sda_i <= '0';
                when 4341 => sda_i <= '0';
                when 4342 => sda_i <= '0';
                when 4343 => sda_i <= '0';
                when 4344 => sda_i <= '0';
                when 4345 => sda_i <= '0';
                when 4346 => sda_i <= '0';
                when 4347 => sda_i <= '0';
                when 4348 => sda_i <= '0';
                when 4349 => sda_i <= '0';
                when 4350 => sda_i <= '0';
                when 4351 => sda_i <= '0';
                when 4352 => sda_i <= '0';
                when 4353 => sda_i <= '0';
                when 4354 => sda_i <= '0';
                when 4355 => sda_i <= '0';
                when 4356 => sda_i <= '0';
                when 4357 => sda_i <= '0';
                when 4358 => sda_i <= '0';
                when 4359 => sda_i <= '0';
                when 4360 => sda_i <= '0';
                when 4361 => sda_i <= '0';
                when 4362 => sda_i <= '0';
                when 4363 => sda_i <= '0';
                when 4364 => sda_i <= '0';
                when 4365 => sda_i <= '0';
                when 4366 => sda_i <= '0';
                when 4367 => sda_i <= '0';
                when 4368 => sda_i <= '0';
                when 4369 => sda_i <= '0';
                when 4370 => sda_i <= '0';
                when 4371 => sda_i <= '0';
                when 4372 => sda_i <= '0';
                when 4373 => sda_i <= '0';
                when 4374 => sda_i <= '0';
                when 4375 => sda_i <= '0';
                when 4376 => sda_i <= '0';
                when 4377 => sda_i <= '0';
                when 4378 => sda_i <= '0';
                when 4379 => sda_i <= '0';
                when 4380 => sda_i <= '0';
                when 4381 => sda_i <= '0';
                when 4382 => sda_i <= '0';
                when 4383 => sda_i <= '0';
                when 4384 => sda_i <= '0';
                when 4385 => sda_i <= '0';
                when 4386 => sda_i <= '0';
                when 4387 => sda_i <= '0';
                when 4388 => sda_i <= '0';
                when 4389 => sda_i <= '0';
                when 4390 => sda_i <= '0';
                when 4391 => sda_i <= '0';
                when 4392 => sda_i <= '0';
                when 4393 => sda_i <= '0';
                when 4394 => sda_i <= '0';
                when 4395 => sda_i <= '0';
                when 4396 => sda_i <= '0';
                when 4397 => sda_i <= '0';
                when 4398 => sda_i <= '0';
                when 4399 => sda_i <= '0';
                when 4400 => sda_i <= '0';
                when 4401 => sda_i <= '0';
                when 4402 => sda_i <= '0';
                when 4403 => sda_i <= '0';
                when 4404 => sda_i <= '0';
                when 4405 => sda_i <= '0';
                when 4406 => sda_i <= '0';
                when 4407 => sda_i <= '0';
                when 4408 => sda_i <= '0';
                when 4409 => sda_i <= '0';
                when 4410 => sda_i <= '0';
                when 4411 => sda_i <= '0';
                when 4412 => sda_i <= '0';
                when 4413 => sda_i <= '0';
                when 4414 => sda_i <= '0';
                when 4415 => sda_i <= '0';
                when 4416 => sda_i <= '0';
                when 4417 => sda_i <= '0';
                when 4418 => sda_i <= '0';
                when 4419 => sda_i <= '0';
                when 4420 => sda_i <= '0';
                when 4421 => sda_i <= '0';
                when 4422 => sda_i <= '0';
                when 4423 => sda_i <= '0';
                when 4424 => sda_i <= '0';
                when 4425 => sda_i <= '0';
                when 4426 => sda_i <= '1';
                when 4427 => sda_i <= '1';
                when 4428 => sda_i <= '0';
                when 4429 => sda_i <= '0';
                when 4430 => sda_i <= '0';
                when 4431 => sda_i <= '0';
                when 4432 => sda_i <= '0';
                when 4433 => sda_i <= '0';
                when 4434 => sda_i <= '0';
                when 4435 => sda_i <= '0';
                when 4436 => sda_i <= '0';
                when 4437 => sda_i <= '0';
                when 4438 => sda_i <= '0';
                when 4439 => sda_i <= '0';
                when 4440 => sda_i <= '0';
                when 4441 => sda_i <= '0';
                when 4442 => sda_i <= '0';
                when 4443 => sda_i <= '0';
                when 4444 => sda_i <= '0';
                when 4445 => sda_i <= '0';
                when 4446 => sda_i <= '0';
                when 4447 => sda_i <= '0';
                when 4448 => sda_i <= '0';
                when 4449 => sda_i <= '0';
                when 4450 => sda_i <= '1';
                when 4451 => sda_i <= '1';
                when 4452 => sda_i <= '1';
                when 4453 => sda_i <= '1';
                when 4454 => sda_i <= '1';
                when 4455 => sda_i <= '1';
                when 4456 => sda_i <= '1';
                when 4457 => sda_i <= '1';
                when 4458 => sda_i <= '1';
                when 4459 => sda_i <= '1';
                when 4460 => sda_i <= '1';
                when 4461 => sda_i <= '0';
                when 4462 => sda_i <= '0';
                when 4463 => sda_i <= '0';
                when 4464 => sda_i <= '0';
                when 4465 => sda_i <= '0';
                when 4466 => sda_i <= '0';
                when 4467 => sda_i <= '0';
                when 4468 => sda_i <= '0';
                when 4469 => sda_i <= '0';
                when 4470 => sda_i <= '0';
                when 4471 => sda_i <= '0';
                when 4472 => sda_i <= '0';
                when 4473 => sda_i <= '0';
                when 4474 => sda_i <= '0';
                when 4475 => sda_i <= '0';
                when 4476 => sda_i <= '0';
                when 4477 => sda_i <= '0';
                when 4478 => sda_i <= '0';
                when 4479 => sda_i <= '0';
                when 4480 => sda_i <= '0';
                when 4481 => sda_i <= '0';
                when 4482 => sda_i <= '0';
                when 4483 => sda_i <= '0';
                when 4484 => sda_i <= '0';
                when 4485 => sda_i <= '0';
                when 4486 => sda_i <= '1';
                when 4487 => sda_i <= '1';
                when 4488 => sda_i <= '1';
                when 4489 => sda_i <= '1';
                when 4490 => sda_i <= '1';
                when 4491 => sda_i <= '1';
                when 4492 => sda_i <= '1';
                when 4493 => sda_i <= '1';
                when 4494 => sda_i <= '1';
                when 4495 => sda_i <= '1';
                when 4496 => sda_i <= '1';
                when 4497 => sda_i <= '0';
                when 4498 => sda_i <= '0';
                when 4499 => sda_i <= '0';
                when 4500 => sda_i <= '0';
                when 4501 => sda_i <= '0';
                when 4502 => sda_i <= '0';
                when 4503 => sda_i <= '0';
                when 4504 => sda_i <= '0';
                when 4505 => sda_i <= '0';
                when 4506 => sda_i <= '0';
                when 4507 => sda_i <= '0';
                when 4508 => sda_i <= '0';
                when 4509 => sda_i <= '0';
                when 4510 => sda_i <= '1';
                when 4511 => sda_i <= '1';
                when 4512 => sda_i <= '1';
                when 4513 => sda_i <= '1';
                when 4514 => sda_i <= '1';
                when 4515 => sda_i <= '1';
                when 4516 => sda_i <= '1';
                when 4517 => sda_i <= '1';
                when 4518 => sda_i <= '1';
                when 4519 => sda_i <= '1';
                when 4520 => sda_i <= '1';
                when 4521 => sda_i <= '0';
                when 4522 => sda_i <= '0';
                when 4523 => sda_i <= '0';
                when 4524 => sda_i <= '0';
                when 4525 => sda_i <= '0';
                when 4526 => sda_i <= '0';
                when 4527 => sda_i <= '0';
                when 4528 => sda_i <= '0';
                when 4529 => sda_i <= '0';
                when 4530 => sda_i <= '0';
                when 4531 => sda_i <= '0';
                when 4532 => sda_i <= '0';
                when 4533 => sda_i <= '0';
                when 4534 => sda_i <= '1';
                when 4535 => sda_i <= '1';
                when 4536 => sda_i <= '0';
                when 4537 => sda_i <= '0';
                when 4538 => sda_i <= '0';
                when 4539 => sda_i <= '0';
                when 4540 => sda_i <= '0';
                when 4541 => sda_i <= '0';
                when 4542 => sda_i <= '0';
                when 4543 => sda_i <= '0';
                when 4544 => sda_i <= '0';
                when 4545 => sda_i <= '0';
                when 4546 => sda_i <= '0';
                when 4547 => sda_i <= '0';
                when 4548 => sda_i <= '0';
                when 4549 => sda_i <= '0';
                when 4550 => sda_i <= '0';
                when 4551 => sda_i <= '0';
                when 4552 => sda_i <= '0';
                when 4553 => sda_i <= '0';
                when 4554 => sda_i <= '0';
                when 4555 => sda_i <= '0';
                when 4556 => sda_i <= '0';
                when 4557 => sda_i <= '0';
                when 4558 => sda_i <= '0';
                when 4559 => sda_i <= '0';
                when 4560 => sda_i <= '0';
                when 4561 => sda_i <= '0';
                when 4562 => sda_i <= '0';
                when 4563 => sda_i <= '0';
                when 4564 => sda_i <= '0';
                when 4565 => sda_i <= '0';
                when 4566 => sda_i <= '0';
                when 4567 => sda_i <= '0';
                when 4568 => sda_i <= '0';
                when 4569 => sda_i <= '0';
                when 4570 => sda_i <= '0';
                when 4571 => sda_i <= '0';
                when 4572 => sda_i <= '0';
                when 4573 => sda_i <= '0';
                when 4574 => sda_i <= '0';
                when 4575 => sda_i <= '0';
                when 4576 => sda_i <= '0';
                when 4577 => sda_i <= '0';
                when 4578 => sda_i <= '0';
                when 4579 => sda_i <= '0';
                when 4580 => sda_i <= '0';
                when 4581 => sda_i <= '0';
                when 4582 => sda_i <= '0';
                when 4583 => sda_i <= '0';
                when 4584 => sda_i <= '0';
                when 4585 => sda_i <= '0';
                when 4586 => sda_i <= '0';
                when 4587 => sda_i <= '0';
                when 4588 => sda_i <= '0';
                when 4589 => sda_i <= '0';
                when 4590 => sda_i <= '0';
                when 4591 => sda_i <= '0';
                when 4592 => sda_i <= '0';
                when 4593 => sda_i <= '0';
                when 4594 => sda_i <= '0';
                when 4595 => sda_i <= '0';
                when 4596 => sda_i <= '0';
                when 4597 => sda_i <= '0';
                when 4598 => sda_i <= '0';
                when 4599 => sda_i <= '0';
                when 4600 => sda_i <= '0';
                when 4601 => sda_i <= '0';
                when 4602 => sda_i <= '0';
                when 4603 => sda_i <= '0';
                when 4604 => sda_i <= '0';
                when 4605 => sda_i <= '0';
                when 4606 => sda_i <= '0';
                when 4607 => sda_i <= '0';
                when 4608 => sda_i <= '0';
                when 4609 => sda_i <= '0';
                when 4610 => sda_i <= '0';
                when 4611 => sda_i <= '0';
                when 4612 => sda_i <= '0';
                when 4613 => sda_i <= '0';
                when 4614 => sda_i <= '0';
                when 4615 => sda_i <= '0';
                when 4616 => sda_i <= '0';
                when 4617 => sda_i <= '0';
                when 4618 => sda_i <= '0';
                when 4619 => sda_i <= '0';
                when 4620 => sda_i <= '0';
                when 4621 => sda_i <= '0';
                when 4622 => sda_i <= '0';
                when 4623 => sda_i <= '0';
                when 4624 => sda_i <= '0';
                when 4625 => sda_i <= '0';
                when 4626 => sda_i <= '0';
                when 4627 => sda_i <= '0';
                when 4628 => sda_i <= '0';
                when 4629 => sda_i <= '0';
                when 4630 => sda_i <= '0';
                when 4631 => sda_i <= '0';
                when 4632 => sda_i <= '0';
                when 4633 => sda_i <= '0';
                when 4634 => sda_i <= '0';
                when 4635 => sda_i <= '0';
                when 4636 => sda_i <= '0';
                when 4637 => sda_i <= '0';
                when 4638 => sda_i <= '0';
                when 4639 => sda_i <= '0';
                when 4640 => sda_i <= '0';
                when 4641 => sda_i <= '0';
                when 4642 => sda_i <= '1';
                when 4643 => sda_i <= '1';
                when 4644 => sda_i <= '0';
                when 4645 => sda_i <= '0';
                when 4646 => sda_i <= '0';
                when 4647 => sda_i <= '0';
                when 4648 => sda_i <= '0';
                when 4649 => sda_i <= '0';
                when 4650 => sda_i <= '0';
                when 4651 => sda_i <= '0';
                when 4652 => sda_i <= '0';
                when 4653 => sda_i <= '0';
                when 4654 => sda_i <= '0';
                when 4655 => sda_i <= '0';
                when 4656 => sda_i <= '0';
                when 4657 => sda_i <= '0';
                when 4658 => sda_i <= '0';
                when 4659 => sda_i <= '0';
                when 4660 => sda_i <= '0';
                when 4661 => sda_i <= '0';
                when 4662 => sda_i <= '0';
                when 4663 => sda_i <= '0';
                when 4664 => sda_i <= '0';
                when 4665 => sda_i <= '0';
                when 4666 => sda_i <= '0';
                when 4667 => sda_i <= '0';
                when 4668 => sda_i <= '0';
                when 4669 => sda_i <= '0';
                when 4670 => sda_i <= '0';
                when 4671 => sda_i <= '0';
                when 4672 => sda_i <= '0';
                when 4673 => sda_i <= '0';
                when 4674 => sda_i <= '0';
                when 4675 => sda_i <= '0';
                when 4676 => sda_i <= '0';
                when 4677 => sda_i <= '0';
                when 4678 => sda_i <= '0';
                when 4679 => sda_i <= '0';
                when 4680 => sda_i <= '0';
                when 4681 => sda_i <= '0';
                when 4682 => sda_i <= '0';
                when 4683 => sda_i <= '0';
                when 4684 => sda_i <= '0';
                when 4685 => sda_i <= '0';
                when 4686 => sda_i <= '0';
                when 4687 => sda_i <= '0';
                when 4688 => sda_i <= '0';
                when 4689 => sda_i <= '0';
                when 4690 => sda_i <= '0';
                when 4691 => sda_i <= '0';
                when 4692 => sda_i <= '0';
                when 4693 => sda_i <= '0';
                when 4694 => sda_i <= '0';
                when 4695 => sda_i <= '0';
                when 4696 => sda_i <= '0';
                when 4697 => sda_i <= '0';
                when 4698 => sda_i <= '0';
                when 4699 => sda_i <= '0';
                when 4700 => sda_i <= '0';
                when 4701 => sda_i <= '0';
                when 4702 => sda_i <= '0';
                when 4703 => sda_i <= '0';
                when 4704 => sda_i <= '0';
                when 4705 => sda_i <= '0';
                when 4706 => sda_i <= '0';
                when 4707 => sda_i <= '0';
                when 4708 => sda_i <= '0';
                when 4709 => sda_i <= '0';
                when 4710 => sda_i <= '0';
                when 4711 => sda_i <= '0';
                when 4712 => sda_i <= '0';
                when 4713 => sda_i <= '0';
                when 4714 => sda_i <= '0';
                when 4715 => sda_i <= '0';
                when 4716 => sda_i <= '0';
                when 4717 => sda_i <= '0';
                when 4718 => sda_i <= '0';
                when 4719 => sda_i <= '0';
                when 4720 => sda_i <= '0';
                when 4721 => sda_i <= '0';
                when 4722 => sda_i <= '0';
                when 4723 => sda_i <= '0';
                when 4724 => sda_i <= '0';
                when 4725 => sda_i <= '0';
                when 4726 => sda_i <= '0';
                when 4727 => sda_i <= '0';
                when 4728 => sda_i <= '0';
                when 4729 => sda_i <= '0';
                when 4730 => sda_i <= '0';
                when 4731 => sda_i <= '0';
                when 4732 => sda_i <= '0';
                when 4733 => sda_i <= '0';
                when 4734 => sda_i <= '0';
                when 4735 => sda_i <= '0';
                when 4736 => sda_i <= '0';
                when 4737 => sda_i <= '0';
                when 4738 => sda_i <= '0';
                when 4739 => sda_i <= '0';
                when 4740 => sda_i <= '0';
                when 4741 => sda_i <= '0';
                when 4742 => sda_i <= '0';
                when 4743 => sda_i <= '0';
                when 4744 => sda_i <= '0';
                when 4745 => sda_i <= '0';
                when 4746 => sda_i <= '0';
                when 4747 => sda_i <= '0';
                when 4748 => sda_i <= '0';
                when 4749 => sda_i <= '0';
                when 4750 => sda_i <= '1';
                when 4751 => sda_i <= '1';
                when 4752 => sda_i <= '0';
                when 4753 => sda_i <= '0';
                when 4754 => sda_i <= '0';
                when 4755 => sda_i <= '0';
                when 4756 => sda_i <= '0';
                when 4757 => sda_i <= '0';
                when 4758 => sda_i <= '0';
                when 4759 => sda_i <= '0';
                when 4760 => sda_i <= '0';
                when 4761 => sda_i <= '0';
                when 4762 => sda_i <= '0';
                when 4763 => sda_i <= '0';
                when 4764 => sda_i <= '0';
                when 4765 => sda_i <= '0';
                when 4766 => sda_i <= '0';
                when 4767 => sda_i <= '0';
                when 4768 => sda_i <= '0';
                when 4769 => sda_i <= '0';
                when 4770 => sda_i <= '0';
                when 4771 => sda_i <= '0';
                when 4772 => sda_i <= '0';
                when 4773 => sda_i <= '0';
                when 4774 => sda_i <= '0';
                when 4775 => sda_i <= '0';
                when 4776 => sda_i <= '0';
                when 4777 => sda_i <= '0';
                when 4778 => sda_i <= '0';
                when 4779 => sda_i <= '0';
                when 4780 => sda_i <= '0';
                when 4781 => sda_i <= '0';
                when 4782 => sda_i <= '0';
                when 4783 => sda_i <= '0';
                when 4784 => sda_i <= '0';
                when 4785 => sda_i <= '0';
                when 4786 => sda_i <= '0';
                when 4787 => sda_i <= '0';
                when 4788 => sda_i <= '0';
                when 4789 => sda_i <= '0';
                when 4790 => sda_i <= '0';
                when 4791 => sda_i <= '0';
                when 4792 => sda_i <= '0';
                when 4793 => sda_i <= '0';
                when 4794 => sda_i <= '0';
                when 4795 => sda_i <= '0';
                when 4796 => sda_i <= '0';
                when 4797 => sda_i <= '0';
                when 4798 => sda_i <= '1';
                when 4799 => sda_i <= '1';
                when 4800 => sda_i <= '1';
                when 4801 => sda_i <= '1';
                when 4802 => sda_i <= '1';
                when 4803 => sda_i <= '1';
                when 4804 => sda_i <= '1';
                when 4805 => sda_i <= '1';
                when 4806 => sda_i <= '1';
                when 4807 => sda_i <= '1';
                when 4808 => sda_i <= '1';
                when 4809 => sda_i <= '0';
                when 4810 => sda_i <= '0';
                when 4811 => sda_i <= '0';
                when 4812 => sda_i <= '0';
                when 4813 => sda_i <= '0';
                when 4814 => sda_i <= '0';
                when 4815 => sda_i <= '0';
                when 4816 => sda_i <= '0';
                when 4817 => sda_i <= '0';
                when 4818 => sda_i <= '0';
                when 4819 => sda_i <= '0';
                when 4820 => sda_i <= '0';
                when 4821 => sda_i <= '0';
                when 4822 => sda_i <= '0';
                when 4823 => sda_i <= '0';
                when 4824 => sda_i <= '0';
                when 4825 => sda_i <= '0';
                when 4826 => sda_i <= '0';
                when 4827 => sda_i <= '0';
                when 4828 => sda_i <= '0';
                when 4829 => sda_i <= '0';
                when 4830 => sda_i <= '0';
                when 4831 => sda_i <= '0';
                when 4832 => sda_i <= '0';
                when 4833 => sda_i <= '0';
                when 4834 => sda_i <= '0';
                when 4835 => sda_i <= '0';
                when 4836 => sda_i <= '0';
                when 4837 => sda_i <= '0';
                when 4838 => sda_i <= '0';
                when 4839 => sda_i <= '0';
                when 4840 => sda_i <= '0';
                when 4841 => sda_i <= '0';
                when 4842 => sda_i <= '0';
                when 4843 => sda_i <= '0';
                when 4844 => sda_i <= '0';
                when 4845 => sda_i <= '0';
                when 4846 => sda_i <= '0';
                when 4847 => sda_i <= '0';
                when 4848 => sda_i <= '0';
                when 4849 => sda_i <= '0';
                when 4850 => sda_i <= '0';
                when 4851 => sda_i <= '0';
                when 4852 => sda_i <= '0';
                when 4853 => sda_i <= '0';
                when 4854 => sda_i <= '0';
                when 4855 => sda_i <= '0';
                when 4856 => sda_i <= '0';
                when 4857 => sda_i <= '0';
                when 4858 => sda_i <= '1';
                when 4859 => sda_i <= '1';
                when 4860 => sda_i <= '0';
                when 4861 => sda_i <= '0';
                when 4862 => sda_i <= '0';
                when 4863 => sda_i <= '0';
                when 4864 => sda_i <= '0';
                when 4865 => sda_i <= '0';
                when 4866 => sda_i <= '0';
                when 4867 => sda_i <= '0';
                when 4868 => sda_i <= '0';
                when 4869 => sda_i <= '0';
                when 4870 => sda_i <= '0';
                when 4871 => sda_i <= '0';
                when 4872 => sda_i <= '0';
                when 4873 => sda_i <= '0';
                when 4874 => sda_i <= '0';
                when 4875 => sda_i <= '0';
                when 4876 => sda_i <= '0';
                when 4877 => sda_i <= '0';
                when 4878 => sda_i <= '0';
                when 4879 => sda_i <= '0';
                when 4880 => sda_i <= '0';
                when 4881 => sda_i <= '0';
                when 4882 => sda_i <= '0';
                when 4883 => sda_i <= '0';
                when 4884 => sda_i <= '0';
                when 4885 => sda_i <= '0';
                when 4886 => sda_i <= '0';
                when 4887 => sda_i <= '0';
                when 4888 => sda_i <= '0';
                when 4889 => sda_i <= '0';
                when 4890 => sda_i <= '0';
                when 4891 => sda_i <= '0';
                when 4892 => sda_i <= '0';
                when 4893 => sda_i <= '0';
                when 4894 => sda_i <= '0';
                when 4895 => sda_i <= '0';
                when 4896 => sda_i <= '0';
                when 4897 => sda_i <= '0';
                when 4898 => sda_i <= '0';
                when 4899 => sda_i <= '0';
                when 4900 => sda_i <= '0';
                when 4901 => sda_i <= '0';
                when 4902 => sda_i <= '0';
                when 4903 => sda_i <= '0';
                when 4904 => sda_i <= '0';
                when 4905 => sda_i <= '0';
                when 4906 => sda_i <= '0';
                when 4907 => sda_i <= '0';
                when 4908 => sda_i <= '0';
                when 4909 => sda_i <= '0';
                when 4910 => sda_i <= '0';
                when 4911 => sda_i <= '0';
                when 4912 => sda_i <= '0';
                when 4913 => sda_i <= '0';
                when 4914 => sda_i <= '0';
                when 4915 => sda_i <= '0';
                when 4916 => sda_i <= '0';
                when 4917 => sda_i <= '0';
                when 4918 => sda_i <= '0';
                when 4919 => sda_i <= '0';
                when 4920 => sda_i <= '0';
                when 4921 => sda_i <= '0';
                when 4922 => sda_i <= '0';
                when 4923 => sda_i <= '0';
                when 4924 => sda_i <= '0';
                when 4925 => sda_i <= '0';
                when 4926 => sda_i <= '0';
                when 4927 => sda_i <= '0';
                when 4928 => sda_i <= '0';
                when 4929 => sda_i <= '0';
                when 4930 => sda_i <= '0';
                when 4931 => sda_i <= '0';
                when 4932 => sda_i <= '0';
                when 4933 => sda_i <= '0';
                when 4934 => sda_i <= '0';
                when 4935 => sda_i <= '0';
                when 4936 => sda_i <= '0';
                when 4937 => sda_i <= '0';
                when 4938 => sda_i <= '0';
                when 4939 => sda_i <= '0';
                when 4940 => sda_i <= '0';
                when 4941 => sda_i <= '0';
                when 4942 => sda_i <= '0';
                when 4943 => sda_i <= '0';
                when 4944 => sda_i <= '0';
                when 4945 => sda_i <= '0';
                when 4946 => sda_i <= '0';
                when 4947 => sda_i <= '0';
                when 4948 => sda_i <= '0';
                when 4949 => sda_i <= '0';
                when 4950 => sda_i <= '0';
                when 4951 => sda_i <= '0';
                when 4952 => sda_i <= '0';
                when 4953 => sda_i <= '0';
                when 4954 => sda_i <= '0';
                when 4955 => sda_i <= '0';
                when 4956 => sda_i <= '0';
                when 4957 => sda_i <= '0';
                when 4958 => sda_i <= '0';
                when 4959 => sda_i <= '0';
                when 4960 => sda_i <= '0';
                when 4961 => sda_i <= '0';
                when 4962 => sda_i <= '0';
                when 4963 => sda_i <= '0';
                when 4964 => sda_i <= '0';
                when 4965 => sda_i <= '0';
                when 4966 => sda_i <= '1';
                when 4967 => sda_i <= '1';
                when 4968 => sda_i <= '0';
                when 4969 => sda_i <= '0';
                when 4970 => sda_i <= '0';
                when 4971 => sda_i <= '0';
                when 4972 => sda_i <= '0';
                when 4973 => sda_i <= '0';
                when 4974 => sda_i <= '0';
                when 4975 => sda_i <= '0';
                when 4976 => sda_i <= '0';
                when 4977 => sda_i <= '0';
                when 4978 => sda_i <= '0';
                when 4979 => sda_i <= '0';
                when 4980 => sda_i <= '0';
                when 4981 => sda_i <= '0';
                when 4982 => sda_i <= '0';
                when 4983 => sda_i <= '0';
                when 4984 => sda_i <= '0';
                when 4985 => sda_i <= '0';
                when 4986 => sda_i <= '0';
                when 4987 => sda_i <= '0';
                when 4988 => sda_i <= '0';
                when 4989 => sda_i <= '0';
                when 4990 => sda_i <= '0';
                when 4991 => sda_i <= '0';
                when 4992 => sda_i <= '0';
                when 4993 => sda_i <= '0';
                when 4994 => sda_i <= '0';
                when 4995 => sda_i <= '0';
                when 4996 => sda_i <= '0';
                when 4997 => sda_i <= '0';
                when 4998 => sda_i <= '0';
                when 4999 => sda_i <= '0';
                when 5000 => sda_i <= '0';
                when 5001 => sda_i <= '0';
                when 5002 => sda_i <= '0';
                when 5003 => sda_i <= '0';
                when 5004 => sda_i <= '0';
                when 5005 => sda_i <= '0';
                when 5006 => sda_i <= '0';
                when 5007 => sda_i <= '0';
                when 5008 => sda_i <= '0';
                when 5009 => sda_i <= '0';
                when 5010 => sda_i <= '0';
                when 5011 => sda_i <= '0';
                when 5012 => sda_i <= '0';
                when 5013 => sda_i <= '0';
                when 5014 => sda_i <= '0';
                when 5015 => sda_i <= '0';
                when 5016 => sda_i <= '0';
                when 5017 => sda_i <= '0';
                when 5018 => sda_i <= '0';
                when 5019 => sda_i <= '0';
                when 5020 => sda_i <= '0';
                when 5021 => sda_i <= '0';
                when 5022 => sda_i <= '0';
                when 5023 => sda_i <= '0';
                when 5024 => sda_i <= '0';
                when 5025 => sda_i <= '0';
                when 5026 => sda_i <= '0';
                when 5027 => sda_i <= '0';
                when 5028 => sda_i <= '0';
                when 5029 => sda_i <= '0';
                when 5030 => sda_i <= '0';
                when 5031 => sda_i <= '0';
                when 5032 => sda_i <= '0';
                when 5033 => sda_i <= '0';
                when 5034 => sda_i <= '0';
                when 5035 => sda_i <= '0';
                when 5036 => sda_i <= '0';
                when 5037 => sda_i <= '0';
                when 5038 => sda_i <= '0';
                when 5039 => sda_i <= '0';
                when 5040 => sda_i <= '0';
                when 5041 => sda_i <= '0';
                when 5042 => sda_i <= '0';
                when 5043 => sda_i <= '0';
                when 5044 => sda_i <= '0';
                when 5045 => sda_i <= '0';
                when 5046 => sda_i <= '0';
                when 5047 => sda_i <= '0';
                when 5048 => sda_i <= '0';
                when 5049 => sda_i <= '0';
                when 5050 => sda_i <= '0';
                when 5051 => sda_i <= '0';
                when 5052 => sda_i <= '0';
                when 5053 => sda_i <= '0';
                when 5054 => sda_i <= '0';
                when 5055 => sda_i <= '0';
                when 5056 => sda_i <= '0';
                when 5057 => sda_i <= '0';
                when 5058 => sda_i <= '0';
                when 5059 => sda_i <= '0';
                when 5060 => sda_i <= '0';
                when 5061 => sda_i <= '0';
                when 5062 => sda_i <= '0';
                when 5063 => sda_i <= '0';
                when 5064 => sda_i <= '0';
                when 5065 => sda_i <= '0';
                when 5066 => sda_i <= '0';
                when 5067 => sda_i <= '0';
                when 5068 => sda_i <= '0';
                when 5069 => sda_i <= '0';
                when 5070 => sda_i <= '0';
                when 5071 => sda_i <= '0';
                when 5072 => sda_i <= '0';
                when 5073 => sda_i <= '0';
                when 5074 => sda_i <= '1';
                when 5075 => sda_i <= '1';
                when 5076 => sda_i <= '0';
                when 5077 => sda_i <= '0';
                when 5078 => sda_i <= '0';
                when 5079 => sda_i <= '0';
                when 5080 => sda_i <= '0';
                when 5081 => sda_i <= '0';
                when 5082 => sda_i <= '0';
                when 5083 => sda_i <= '0';
                when 5084 => sda_i <= '0';
                when 5085 => sda_i <= '0';
                when 5086 => sda_i <= '0';
                when 5087 => sda_i <= '0';
                when 5088 => sda_i <= '0';
                when 5089 => sda_i <= '0';
                when 5090 => sda_i <= '0';
                when 5091 => sda_i <= '0';
                when 5092 => sda_i <= '0';
                when 5093 => sda_i <= '0';
                when 5094 => sda_i <= '0';
                when 5095 => sda_i <= '0';
                when 5096 => sda_i <= '0';
                when 5097 => sda_i <= '0';
                when 5098 => sda_i <= '0';
                when 5099 => sda_i <= '0';
                when 5100 => sda_i <= '0';
                when 5101 => sda_i <= '0';
                when 5102 => sda_i <= '0';
                when 5103 => sda_i <= '0';
                when 5104 => sda_i <= '0';
                when 5105 => sda_i <= '0';
                when 5106 => sda_i <= '0';
                when 5107 => sda_i <= '0';
                when 5108 => sda_i <= '0';
                when 5109 => sda_i <= '0';
                when 5110 => sda_i <= '0';
                when 5111 => sda_i <= '0';
                when 5112 => sda_i <= '0';
                when 5113 => sda_i <= '0';
                when 5114 => sda_i <= '0';
                when 5115 => sda_i <= '0';
                when 5116 => sda_i <= '0';
                when 5117 => sda_i <= '0';
                when 5118 => sda_i <= '0';
                when 5119 => sda_i <= '0';
                when 5120 => sda_i <= '0';
                when 5121 => sda_i <= '0';
                when 5122 => sda_i <= '0';
                when 5123 => sda_i <= '0';
                when 5124 => sda_i <= '0';
                when 5125 => sda_i <= '0';
                when 5126 => sda_i <= '0';
                when 5127 => sda_i <= '0';
                when 5128 => sda_i <= '0';
                when 5129 => sda_i <= '0';
                when 5130 => sda_i <= '0';
                when 5131 => sda_i <= '0';
                when 5132 => sda_i <= '0';
                when 5133 => sda_i <= '0';
                when 5134 => sda_i <= '0';
                when 5135 => sda_i <= '0';
                when 5136 => sda_i <= '0';
                when 5137 => sda_i <= '0';
                when 5138 => sda_i <= '0';
                when 5139 => sda_i <= '0';
                when 5140 => sda_i <= '0';
                when 5141 => sda_i <= '0';
                when 5142 => sda_i <= '0';
                when 5143 => sda_i <= '0';
                when 5144 => sda_i <= '0';
                when 5145 => sda_i <= '0';
                when 5146 => sda_i <= '0';
                when 5147 => sda_i <= '0';
                when 5148 => sda_i <= '0';
                when 5149 => sda_i <= '0';
                when 5150 => sda_i <= '0';
                when 5151 => sda_i <= '0';
                when 5152 => sda_i <= '0';
                when 5153 => sda_i <= '0';
                when 5154 => sda_i <= '0';
                when 5155 => sda_i <= '0';
                when 5156 => sda_i <= '0';
                when 5157 => sda_i <= '0';
                when 5158 => sda_i <= '0';
                when 5159 => sda_i <= '0';
                when 5160 => sda_i <= '0';
                when 5161 => sda_i <= '0';
                when 5162 => sda_i <= '0';
                when 5163 => sda_i <= '0';
                when 5164 => sda_i <= '0';
                when 5165 => sda_i <= '0';
                when 5166 => sda_i <= '0';
                when 5167 => sda_i <= '0';
                when 5168 => sda_i <= '0';
                when 5169 => sda_i <= '0';
                when 5170 => sda_i <= '0';
                when 5171 => sda_i <= '0';
                when 5172 => sda_i <= '0';
                when 5173 => sda_i <= '0';
                when 5174 => sda_i <= '0';
                when 5175 => sda_i <= '0';
                when 5176 => sda_i <= '0';
                when 5177 => sda_i <= '0';
                when 5178 => sda_i <= '0';
                when 5179 => sda_i <= '0';
                when 5180 => sda_i <= '0';
                when 5181 => sda_i <= '0';
                when 5182 => sda_i <= '1';
                when 5183 => sda_i <= '1';
                when 5184 => sda_i <= '0';
                when 5185 => sda_i <= '0';
                when 5186 => sda_i <= '0';
                when 5187 => sda_i <= '0';
                when 5188 => sda_i <= '0';
                when 5189 => sda_i <= '0';
                when 5190 => sda_i <= '0';
                when 5191 => sda_i <= '0';
                when 5192 => sda_i <= '0';
                when 5193 => sda_i <= '0';
                when 5194 => sda_i <= '0';
                when 5195 => sda_i <= '0';
                when 5196 => sda_i <= '0';
                when 5197 => sda_i <= '0';
                when 5198 => sda_i <= '0';
                when 5199 => sda_i <= '0';
                when 5200 => sda_i <= '0';
                when 5201 => sda_i <= '0';
                when 5202 => sda_i <= '0';
                when 5203 => sda_i <= '0';
                when 5204 => sda_i <= '0';
                when 5205 => sda_i <= '0';
                when 5206 => sda_i <= '0';
                when 5207 => sda_i <= '0';
                when 5208 => sda_i <= '0';
                when 5209 => sda_i <= '0';
                when 5210 => sda_i <= '0';
                when 5211 => sda_i <= '0';
                when 5212 => sda_i <= '0';
                when 5213 => sda_i <= '0';
                when 5214 => sda_i <= '0';
                when 5215 => sda_i <= '0';
                when 5216 => sda_i <= '0';
                when 5217 => sda_i <= '0';
                when 5218 => sda_i <= '0';
                when 5219 => sda_i <= '0';
                when 5220 => sda_i <= '0';
                when 5221 => sda_i <= '0';
                when 5222 => sda_i <= '0';
                when 5223 => sda_i <= '0';
                when 5224 => sda_i <= '0';
                when 5225 => sda_i <= '0';
                when 5226 => sda_i <= '0';
                when 5227 => sda_i <= '0';
                when 5228 => sda_i <= '0';
                when 5229 => sda_i <= '0';
                when 5230 => sda_i <= '0';
                when 5231 => sda_i <= '0';
                when 5232 => sda_i <= '0';
                when 5233 => sda_i <= '0';
                when 5234 => sda_i <= '0';
                when 5235 => sda_i <= '0';
                when 5236 => sda_i <= '0';
                when 5237 => sda_i <= '0';
                when 5238 => sda_i <= '0';
                when 5239 => sda_i <= '0';
                when 5240 => sda_i <= '0';
                when 5241 => sda_i <= '0';
                when 5242 => sda_i <= '0';
                when 5243 => sda_i <= '0';
                when 5244 => sda_i <= '0';
                when 5245 => sda_i <= '0';
                when 5246 => sda_i <= '0';
                when 5247 => sda_i <= '0';
                when 5248 => sda_i <= '0';
                when 5249 => sda_i <= '0';
                when 5250 => sda_i <= '0';
                when 5251 => sda_i <= '0';
                when 5252 => sda_i <= '0';
                when 5253 => sda_i <= '0';
                when 5254 => sda_i <= '0';
                when 5255 => sda_i <= '0';
                when 5256 => sda_i <= '0';
                when 5257 => sda_i <= '0';
                when 5258 => sda_i <= '0';
                when 5259 => sda_i <= '0';
                when 5260 => sda_i <= '0';
                when 5261 => sda_i <= '0';
                when 5262 => sda_i <= '0';
                when 5263 => sda_i <= '0';
                when 5264 => sda_i <= '0';
                when 5265 => sda_i <= '0';
                when 5266 => sda_i <= '0';
                when 5267 => sda_i <= '0';
                when 5268 => sda_i <= '0';
                when 5269 => sda_i <= '0';
                when 5270 => sda_i <= '0';
                when 5271 => sda_i <= '0';
                when 5272 => sda_i <= '0';
                when 5273 => sda_i <= '0';
                when 5274 => sda_i <= '0';
                when 5275 => sda_i <= '0';
                when 5276 => sda_i <= '0';
                when 5277 => sda_i <= '0';
                when 5278 => sda_i <= '0';
                when 5279 => sda_i <= '0';
                when 5280 => sda_i <= '0';
                when 5281 => sda_i <= '0';
                when 5282 => sda_i <= '0';
                when 5283 => sda_i <= '0';
                when 5284 => sda_i <= '0';
                when 5285 => sda_i <= '0';
                when 5286 => sda_i <= '0';
                when 5287 => sda_i <= '0';
                when 5288 => sda_i <= '0';
                when 5289 => sda_i <= '0';
                when 5290 => sda_i <= '1';
                when 5291 => sda_i <= '1';
                when 5292 => sda_i <= '0';
                when 5293 => sda_i <= '0';
                when 5294 => sda_i <= '0';
                when 5295 => sda_i <= '0';
                when 5296 => sda_i <= '0';
                when 5297 => sda_i <= '0';
                when 5298 => sda_i <= '0';
                when 5299 => sda_i <= '0';
                when 5300 => sda_i <= '0';
                when 5301 => sda_i <= '0';
                when 5302 => sda_i <= '0';
                when 5303 => sda_i <= '0';
                when 5304 => sda_i <= '0';
                when 5305 => sda_i <= '0';
                when 5306 => sda_i <= '0';
                when 5307 => sda_i <= '0';
                when 5308 => sda_i <= '0';
                when 5309 => sda_i <= '0';
                when 5310 => sda_i <= '0';
                when 5311 => sda_i <= '0';
                when 5312 => sda_i <= '0';
                when 5313 => sda_i <= '0';
                when 5314 => sda_i <= '0';
                when 5315 => sda_i <= '0';
                when 5316 => sda_i <= '0';
                when 5317 => sda_i <= '0';
                when 5318 => sda_i <= '0';
                when 5319 => sda_i <= '0';
                when 5320 => sda_i <= '0';
                when 5321 => sda_i <= '0';
                when 5322 => sda_i <= '0';
                when 5323 => sda_i <= '0';
                when 5324 => sda_i <= '0';
                when 5325 => sda_i <= '0';
                when 5326 => sda_i <= '0';
                when 5327 => sda_i <= '0';
                when 5328 => sda_i <= '0';
                when 5329 => sda_i <= '0';
                when 5330 => sda_i <= '0';
                when 5331 => sda_i <= '0';
                when 5332 => sda_i <= '0';
                when 5333 => sda_i <= '0';
                when 5334 => sda_i <= '0';
                when 5335 => sda_i <= '0';
                when 5336 => sda_i <= '0';
                when 5337 => sda_i <= '0';
                when 5338 => sda_i <= '0';
                when 5339 => sda_i <= '0';
                when 5340 => sda_i <= '0';
                when 5341 => sda_i <= '0';
                when 5342 => sda_i <= '0';
                when 5343 => sda_i <= '0';
                when 5344 => sda_i <= '0';
                when 5345 => sda_i <= '0';
                when 5346 => sda_i <= '0';
                when 5347 => sda_i <= '0';
                when 5348 => sda_i <= '0';
                when 5349 => sda_i <= '0';
                when 5350 => sda_i <= '0';
                when 5351 => sda_i <= '0';
                when 5352 => sda_i <= '0';
                when 5353 => sda_i <= '0';
                when 5354 => sda_i <= '0';
                when 5355 => sda_i <= '0';
                when 5356 => sda_i <= '0';
                when 5357 => sda_i <= '0';
                when 5358 => sda_i <= '0';
                when 5359 => sda_i <= '0';
                when 5360 => sda_i <= '0';
                when 5361 => sda_i <= '0';
                when 5362 => sda_i <= '0';
                when 5363 => sda_i <= '0';
                when 5364 => sda_i <= '0';
                when 5365 => sda_i <= '0';
                when 5366 => sda_i <= '0';
                when 5367 => sda_i <= '0';
                when 5368 => sda_i <= '0';
                when 5369 => sda_i <= '0';
                when 5370 => sda_i <= '0';
                when 5371 => sda_i <= '0';
                when 5372 => sda_i <= '0';
                when 5373 => sda_i <= '0';
                when 5374 => sda_i <= '0';
                when 5375 => sda_i <= '0';
                when 5376 => sda_i <= '0';
                when 5377 => sda_i <= '0';
                when 5378 => sda_i <= '0';
                when 5379 => sda_i <= '0';
                when 5380 => sda_i <= '0';
                when 5381 => sda_i <= '0';
                when 5382 => sda_i <= '0';
                when 5383 => sda_i <= '0';
                when 5384 => sda_i <= '0';
                when 5385 => sda_i <= '0';
                when 5386 => sda_i <= '0';
                when 5387 => sda_i <= '0';
                when 5388 => sda_i <= '0';
                when 5389 => sda_i <= '0';
                when 5390 => sda_i <= '0';
                when 5391 => sda_i <= '0';
                when 5392 => sda_i <= '0';
                when 5393 => sda_i <= '0';
                when 5394 => sda_i <= '0';
                when 5395 => sda_i <= '0';
                when 5396 => sda_i <= '0';
                when 5397 => sda_i <= '0';
                when 5398 => sda_i <= '1';
                when 5399 => sda_i <= '1';
                when 5400 => sda_i <= '0';
                when 5401 => sda_i <= '0';
                when 5402 => sda_i <= '0';
                when 5403 => sda_i <= '0';
                when 5404 => sda_i <= '0';
                when 5405 => sda_i <= '0';
                when 5406 => sda_i <= '0';
                when 5407 => sda_i <= '0';
                when 5408 => sda_i <= '0';
                when 5409 => sda_i <= '0';
                when 5410 => sda_i <= '0';
                when 5411 => sda_i <= '0';
                when 5412 => sda_i <= '0';
                when 5413 => sda_i <= '0';
                when 5414 => sda_i <= '0';
                when 5415 => sda_i <= '0';
                when 5416 => sda_i <= '0';
                when 5417 => sda_i <= '0';
                when 5418 => sda_i <= '0';
                when 5419 => sda_i <= '0';
                when 5420 => sda_i <= '0';
                when 5421 => sda_i <= '0';
                when 5422 => sda_i <= '0';
                when 5423 => sda_i <= '0';
                when 5424 => sda_i <= '0';
                when 5425 => sda_i <= '0';
                when 5426 => sda_i <= '0';
                when 5427 => sda_i <= '0';
                when 5428 => sda_i <= '0';
                when 5429 => sda_i <= '0';
                when 5430 => sda_i <= '0';
                when 5431 => sda_i <= '0';
                when 5432 => sda_i <= '0';
                when 5433 => sda_i <= '0';
                when 5434 => sda_i <= '0';
                when 5435 => sda_i <= '0';
                when 5436 => sda_i <= '0';
                when 5437 => sda_i <= '0';
                when 5438 => sda_i <= '0';
                when 5439 => sda_i <= '0';
                when 5440 => sda_i <= '0';
                when 5441 => sda_i <= '0';
                when 5442 => sda_i <= '0';
                when 5443 => sda_i <= '0';
                when 5444 => sda_i <= '0';
                when 5445 => sda_i <= '0';
                when 5446 => sda_i <= '0';
                when 5447 => sda_i <= '0';
                when 5448 => sda_i <= '0';
                when 5449 => sda_i <= '0';
                when 5450 => sda_i <= '0';
                when 5451 => sda_i <= '0';
                when 5452 => sda_i <= '0';
                when 5453 => sda_i <= '0';
                when 5454 => sda_i <= '0';
                when 5455 => sda_i <= '0';
                when 5456 => sda_i <= '0';
                when 5457 => sda_i <= '0';
                when 5458 => sda_i <= '0';
                when 5459 => sda_i <= '0';
                when 5460 => sda_i <= '0';
                when 5461 => sda_i <= '0';
                when 5462 => sda_i <= '0';
                when 5463 => sda_i <= '0';
                when 5464 => sda_i <= '0';
                when 5465 => sda_i <= '0';
                when 5466 => sda_i <= '0';
                when 5467 => sda_i <= '0';
                when 5468 => sda_i <= '0';
                when 5469 => sda_i <= '0';
                when 5470 => sda_i <= '0';
                when 5471 => sda_i <= '0';
                when 5472 => sda_i <= '0';
                when 5473 => sda_i <= '0';
                when 5474 => sda_i <= '0';
                when 5475 => sda_i <= '0';
                when 5476 => sda_i <= '0';
                when 5477 => sda_i <= '0';
                when 5478 => sda_i <= '0';
                when 5479 => sda_i <= '0';
                when 5480 => sda_i <= '0';
                when 5481 => sda_i <= '0';
                when 5482 => sda_i <= '0';
                when 5483 => sda_i <= '0';
                when 5484 => sda_i <= '0';
                when 5485 => sda_i <= '0';
                when 5486 => sda_i <= '0';
                when 5487 => sda_i <= '0';
                when 5488 => sda_i <= '0';
                when 5489 => sda_i <= '0';
                when 5490 => sda_i <= '0';
                when 5491 => sda_i <= '0';
                when 5492 => sda_i <= '0';
                when 5493 => sda_i <= '0';
                when 5494 => sda_i <= '0';
                when 5495 => sda_i <= '0';
                when 5496 => sda_i <= '0';
                when 5497 => sda_i <= '0';
                when 5498 => sda_i <= '0';
                when 5499 => sda_i <= '0';
                when 5500 => sda_i <= '0';
                when 5501 => sda_i <= '0';
                when 5502 => sda_i <= '0';
                when 5503 => sda_i <= '0';
                when 5504 => sda_i <= '0';
                when 5505 => sda_i <= '0';
                when 5506 => sda_i <= '1';
                when 5507 => sda_i <= '1';
                when 5508 => sda_i <= '0';
                when 5509 => sda_i <= '0';
                when 5510 => sda_i <= '0';
                when 5511 => sda_i <= '0';
                when 5512 => sda_i <= '0';
                when 5513 => sda_i <= '0';
                when 5514 => sda_i <= '0';
                when 5515 => sda_i <= '0';
                when 5516 => sda_i <= '0';
                when 5517 => sda_i <= '0';
                when 5518 => sda_i <= '0';
                when 5519 => sda_i <= '0';
                when 5520 => sda_i <= '0';
                when 5521 => sda_i <= '0';
                when 5522 => sda_i <= '0';
                when 5523 => sda_i <= '0';
                when 5524 => sda_i <= '0';
                when 5525 => sda_i <= '0';
                when 5526 => sda_i <= '0';
                when 5527 => sda_i <= '0';
                when 5528 => sda_i <= '0';
                when 5529 => sda_i <= '0';
                when 5530 => sda_i <= '0';
                when 5531 => sda_i <= '0';
                when 5532 => sda_i <= '0';
                when 5533 => sda_i <= '0';
                when 5534 => sda_i <= '0';
                when 5535 => sda_i <= '0';
                when 5536 => sda_i <= '0';
                when 5537 => sda_i <= '0';
                when 5538 => sda_i <= '0';
                when 5539 => sda_i <= '0';
                when 5540 => sda_i <= '0';
                when 5541 => sda_i <= '0';
                when 5542 => sda_i <= '0';
                when 5543 => sda_i <= '0';
                when 5544 => sda_i <= '0';
                when 5545 => sda_i <= '0';
                when 5546 => sda_i <= '0';
                when 5547 => sda_i <= '0';
                when 5548 => sda_i <= '0';
                when 5549 => sda_i <= '0';
                when 5550 => sda_i <= '0';
                when 5551 => sda_i <= '0';
                when 5552 => sda_i <= '0';
                when 5553 => sda_i <= '0';
                when 5554 => sda_i <= '0';
                when 5555 => sda_i <= '0';
                when 5556 => sda_i <= '0';
                when 5557 => sda_i <= '0';
                when 5558 => sda_i <= '0';
                when 5559 => sda_i <= '0';
                when 5560 => sda_i <= '0';
                when 5561 => sda_i <= '0';
                when 5562 => sda_i <= '0';
                when 5563 => sda_i <= '0';
                when 5564 => sda_i <= '0';
                when 5565 => sda_i <= '0';
                when 5566 => sda_i <= '0';
                when 5567 => sda_i <= '0';
                when 5568 => sda_i <= '0';
                when 5569 => sda_i <= '0';
                when 5570 => sda_i <= '0';
                when 5571 => sda_i <= '0';
                when 5572 => sda_i <= '0';
                when 5573 => sda_i <= '0';
                when 5574 => sda_i <= '0';
                when 5575 => sda_i <= '0';
                when 5576 => sda_i <= '0';
                when 5577 => sda_i <= '0';
                when 5578 => sda_i <= '0';
                when 5579 => sda_i <= '0';
                when 5580 => sda_i <= '0';
                when 5581 => sda_i <= '0';
                when 5582 => sda_i <= '0';
                when 5583 => sda_i <= '0';
                when 5584 => sda_i <= '0';
                when 5585 => sda_i <= '0';
                when 5586 => sda_i <= '0';
                when 5587 => sda_i <= '0';
                when 5588 => sda_i <= '0';
                when 5589 => sda_i <= '0';
                when 5590 => sda_i <= '0';
                when 5591 => sda_i <= '0';
                when 5592 => sda_i <= '0';
                when 5593 => sda_i <= '0';
                when 5594 => sda_i <= '0';
                when 5595 => sda_i <= '0';
                when 5596 => sda_i <= '0';
                when 5597 => sda_i <= '0';
                when 5598 => sda_i <= '0';
                when 5599 => sda_i <= '0';
                when 5600 => sda_i <= '0';
                when 5601 => sda_i <= '0';
                when 5602 => sda_i <= '0';
                when 5603 => sda_i <= '0';
                when 5604 => sda_i <= '0';
                when 5605 => sda_i <= '0';
                when 5606 => sda_i <= '0';
                when 5607 => sda_i <= '0';
                when 5608 => sda_i <= '0';
                when 5609 => sda_i <= '0';
                when 5610 => sda_i <= '0';
                when 5611 => sda_i <= '0';
                when 5612 => sda_i <= '0';
                when 5613 => sda_i <= '0';
                when 5614 => sda_i <= '1';
                when 5615 => sda_i <= '1';
                when 5616 => sda_i <= '0';
                when 5617 => sda_i <= '0';
                when 5618 => sda_i <= '0';
                when 5619 => sda_i <= '0';
                when 5620 => sda_i <= '0';
                when 5621 => sda_i <= '0';
                when 5622 => sda_i <= '0';
                when 5623 => sda_i <= '0';
                when 5624 => sda_i <= '0';
                when 5625 => sda_i <= '0';
                when 5626 => sda_i <= '0';
                when 5627 => sda_i <= '0';
                when 5628 => sda_i <= '0';
                when 5629 => sda_i <= '0';
                when 5630 => sda_i <= '0';
                when 5631 => sda_i <= '0';
                when 5632 => sda_i <= '0';
                when 5633 => sda_i <= '0';
                when 5634 => sda_i <= '0';
                when 5635 => sda_i <= '0';
                when 5636 => sda_i <= '0';
                when 5637 => sda_i <= '0';
                when 5638 => sda_i <= '0';
                when 5639 => sda_i <= '0';
                when 5640 => sda_i <= '0';
                when 5641 => sda_i <= '0';
                when 5642 => sda_i <= '0';
                when 5643 => sda_i <= '0';
                when 5644 => sda_i <= '0';
                when 5645 => sda_i <= '0';
                when 5646 => sda_i <= '0';
                when 5647 => sda_i <= '0';
                when 5648 => sda_i <= '0';
                when 5649 => sda_i <= '0';
                when 5650 => sda_i <= '0';
                when 5651 => sda_i <= '0';
                when 5652 => sda_i <= '0';
                when 5653 => sda_i <= '0';
                when 5654 => sda_i <= '0';
                when 5655 => sda_i <= '0';
                when 5656 => sda_i <= '0';
                when 5657 => sda_i <= '0';
                when 5658 => sda_i <= '0';
                when 5659 => sda_i <= '0';
                when 5660 => sda_i <= '0';
                when 5661 => sda_i <= '0';
                when 5662 => sda_i <= '0';
                when 5663 => sda_i <= '0';
                when 5664 => sda_i <= '0';
                when 5665 => sda_i <= '0';
                when 5666 => sda_i <= '0';
                when 5667 => sda_i <= '0';
                when 5668 => sda_i <= '0';
                when 5669 => sda_i <= '0';
                when 5670 => sda_i <= '0';
                when 5671 => sda_i <= '0';
                when 5672 => sda_i <= '0';
                when 5673 => sda_i <= '0';
                when 5674 => sda_i <= '0';
                when 5675 => sda_i <= '0';
                when 5676 => sda_i <= '0';
                when 5677 => sda_i <= '0';
                when 5678 => sda_i <= '0';
                when 5679 => sda_i <= '0';
                when 5680 => sda_i <= '0';
                when 5681 => sda_i <= '0';
                when 5682 => sda_i <= '0';
                when 5683 => sda_i <= '0';
                when 5684 => sda_i <= '0';
                when 5685 => sda_i <= '0';
                when 5686 => sda_i <= '0';
                when 5687 => sda_i <= '0';
                when 5688 => sda_i <= '0';
                when 5689 => sda_i <= '0';
                when 5690 => sda_i <= '0';
                when 5691 => sda_i <= '0';
                when 5692 => sda_i <= '0';
                when 5693 => sda_i <= '0';
                when 5694 => sda_i <= '0';
                when 5695 => sda_i <= '0';
                when 5696 => sda_i <= '0';
                when 5697 => sda_i <= '0';
                when 5698 => sda_i <= '0';
                when 5699 => sda_i <= '0';
                when 5700 => sda_i <= '0';
                when 5701 => sda_i <= '0';
                when 5702 => sda_i <= '0';
                when 5703 => sda_i <= '0';
                when 5704 => sda_i <= '0';
                when 5705 => sda_i <= '0';
                when 5706 => sda_i <= '0';
                when 5707 => sda_i <= '0';
                when 5708 => sda_i <= '0';
                when 5709 => sda_i <= '0';
                when 5710 => sda_i <= '0';
                when 5711 => sda_i <= '0';
                when 5712 => sda_i <= '0';
                when 5713 => sda_i <= '0';
                when 5714 => sda_i <= '0';
                when 5715 => sda_i <= '0';
                when 5716 => sda_i <= '0';
                when 5717 => sda_i <= '0';
                when 5718 => sda_i <= '0';
                when 5719 => sda_i <= '0';
                when 5720 => sda_i <= '0';
                when 5721 => sda_i <= '0';
                when 5722 => sda_i <= '1';
                when 5723 => sda_i <= '1';
                when 5724 => sda_i <= '0';
                when 5725 => sda_i <= '0';
                when 5726 => sda_i <= '0';
                when 5727 => sda_i <= '0';
                when 5728 => sda_i <= '0';
                when 5729 => sda_i <= '0';
                when 5730 => sda_i <= '0';
                when 5731 => sda_i <= '0';
                when 5732 => sda_i <= '0';
                when 5733 => sda_i <= '0';
                when 5734 => sda_i <= '0';
                when 5735 => sda_i <= '0';
                when 5736 => sda_i <= '0';
                when 5737 => sda_i <= '0';
                when 5738 => sda_i <= '0';
                when 5739 => sda_i <= '0';
                when 5740 => sda_i <= '0';
                when 5741 => sda_i <= '0';
                when 5742 => sda_i <= '0';
                when 5743 => sda_i <= '0';
                when 5744 => sda_i <= '0';
                when 5745 => sda_i <= '0';
                when 5746 => sda_i <= '0';
                when 5747 => sda_i <= '0';
                when 5748 => sda_i <= '0';
                when 5749 => sda_i <= '0';
                when 5750 => sda_i <= '0';
                when 5751 => sda_i <= '0';
                when 5752 => sda_i <= '0';
                when 5753 => sda_i <= '0';
                when 5754 => sda_i <= '0';
                when 5755 => sda_i <= '0';
                when 5756 => sda_i <= '0';
                when 5757 => sda_i <= '0';
                when 5758 => sda_i <= '0';
                when 5759 => sda_i <= '0';
                when 5760 => sda_i <= '0';
                when 5761 => sda_i <= '0';
                when 5762 => sda_i <= '0';
                when 5763 => sda_i <= '0';
                when 5764 => sda_i <= '0';
                when 5765 => sda_i <= '0';
                when 5766 => sda_i <= '0';
                when 5767 => sda_i <= '0';
                when 5768 => sda_i <= '0';
                when 5769 => sda_i <= '0';
                when 5770 => sda_i <= '0';
                when 5771 => sda_i <= '0';
                when 5772 => sda_i <= '0';
                when 5773 => sda_i <= '0';
                when 5774 => sda_i <= '0';
                when 5775 => sda_i <= '0';
                when 5776 => sda_i <= '0';
                when 5777 => sda_i <= '0';
                when 5778 => sda_i <= '0';
                when 5779 => sda_i <= '0';
                when 5780 => sda_i <= '0';
                when 5781 => sda_i <= '0';
                when 5782 => sda_i <= '0';
                when 5783 => sda_i <= '0';
                when 5784 => sda_i <= '0';
                when 5785 => sda_i <= '0';
                when 5786 => sda_i <= '0';
                when 5787 => sda_i <= '0';
                when 5788 => sda_i <= '0';
                when 5789 => sda_i <= '0';
                when 5790 => sda_i <= '0';
                when 5791 => sda_i <= '0';
                when 5792 => sda_i <= '0';
                when 5793 => sda_i <= '0';
                when 5794 => sda_i <= '0';
                when 5795 => sda_i <= '0';
                when 5796 => sda_i <= '0';
                when 5797 => sda_i <= '0';
                when 5798 => sda_i <= '0';
                when 5799 => sda_i <= '0';
                when 5800 => sda_i <= '0';
                when 5801 => sda_i <= '0';
                when 5802 => sda_i <= '0';
                when 5803 => sda_i <= '0';
                when 5804 => sda_i <= '0';
                when 5805 => sda_i <= '0';
                when 5806 => sda_i <= '0';
                when 5807 => sda_i <= '0';
                when 5808 => sda_i <= '0';
                when 5809 => sda_i <= '0';
                when 5810 => sda_i <= '0';
                when 5811 => sda_i <= '0';
                when 5812 => sda_i <= '0';
                when 5813 => sda_i <= '0';
                when 5814 => sda_i <= '0';
                when 5815 => sda_i <= '0';
                when 5816 => sda_i <= '0';
                when 5817 => sda_i <= '0';
                when 5818 => sda_i <= '0';
                when 5819 => sda_i <= '0';
                when 5820 => sda_i <= '0';
                when 5821 => sda_i <= '0';
                when 5822 => sda_i <= '0';
                when 5823 => sda_i <= '0';
                when 5824 => sda_i <= '0';
                when 5825 => sda_i <= '0';
                when 5826 => sda_i <= '0';
                when 5827 => sda_i <= '0';
                when 5828 => sda_i <= '0';
                when 5829 => sda_i <= '0';
                when 5830 => sda_i <= '1';
                when 5831 => sda_i <= '1';
                when 5832 => sda_i <= '0';
                when 5833 => sda_i <= '0';
                when 5834 => sda_i <= '0';
                when 5835 => sda_i <= '0';
                when 5836 => sda_i <= '0';
                when 5837 => sda_i <= '0';
                when 5838 => sda_i <= '0';
                when 5839 => sda_i <= '0';
                when 5840 => sda_i <= '0';
                when 5841 => sda_i <= '0';
                when 5842 => sda_i <= '0';
                when 5843 => sda_i <= '0';
                when 5844 => sda_i <= '0';
                when 5845 => sda_i <= '0';
                when 5846 => sda_i <= '0';
                when 5847 => sda_i <= '0';
                when 5848 => sda_i <= '0';
                when 5849 => sda_i <= '0';
                when 5850 => sda_i <= '0';
                when 5851 => sda_i <= '0';
                when 5852 => sda_i <= '0';
                when 5853 => sda_i <= '0';
                when 5854 => sda_i <= '0';
                when 5855 => sda_i <= '0';
                when 5856 => sda_i <= '0';
                when 5857 => sda_i <= '0';
                when 5858 => sda_i <= '0';
                when 5859 => sda_i <= '0';
                when 5860 => sda_i <= '0';
                when 5861 => sda_i <= '0';
                when 5862 => sda_i <= '0';
                when 5863 => sda_i <= '0';
                when 5864 => sda_i <= '0';
                when 5865 => sda_i <= '0';
                when 5866 => sda_i <= '0';
                when 5867 => sda_i <= '0';
                when 5868 => sda_i <= '0';
                when 5869 => sda_i <= '0';
                when 5870 => sda_i <= '0';
                when 5871 => sda_i <= '0';
                when 5872 => sda_i <= '0';
                when 5873 => sda_i <= '0';
                when 5874 => sda_i <= '0';
                when 5875 => sda_i <= '0';
                when 5876 => sda_i <= '0';
                when 5877 => sda_i <= '0';
                when 5878 => sda_i <= '0';
                when 5879 => sda_i <= '0';
                when 5880 => sda_i <= '0';
                when 5881 => sda_i <= '0';
                when 5882 => sda_i <= '0';
                when 5883 => sda_i <= '0';
                when 5884 => sda_i <= '0';
                when 5885 => sda_i <= '0';
                when 5886 => sda_i <= '0';
                when 5887 => sda_i <= '0';
                when 5888 => sda_i <= '0';
                when 5889 => sda_i <= '0';
                when 5890 => sda_i <= '0';
                when 5891 => sda_i <= '0';
                when 5892 => sda_i <= '0';
                when 5893 => sda_i <= '0';
                when 5894 => sda_i <= '0';
                when 5895 => sda_i <= '0';
                when 5896 => sda_i <= '0';
                when 5897 => sda_i <= '0';
                when 5898 => sda_i <= '0';
                when 5899 => sda_i <= '0';
                when 5900 => sda_i <= '0';
                when 5901 => sda_i <= '0';
                when 5902 => sda_i <= '0';
                when 5903 => sda_i <= '0';
                when 5904 => sda_i <= '0';
                when 5905 => sda_i <= '0';
                when 5906 => sda_i <= '0';
                when 5907 => sda_i <= '0';
                when 5908 => sda_i <= '0';
                when 5909 => sda_i <= '0';
                when 5910 => sda_i <= '0';
                when 5911 => sda_i <= '0';
                when 5912 => sda_i <= '0';
                when 5913 => sda_i <= '0';
                when 5914 => sda_i <= '0';
                when 5915 => sda_i <= '0';
                when 5916 => sda_i <= '0';
                when 5917 => sda_i <= '0';
                when 5918 => sda_i <= '0';
                when 5919 => sda_i <= '0';
                when 5920 => sda_i <= '0';
                when 5921 => sda_i <= '0';
                when 5922 => sda_i <= '0';
                when 5923 => sda_i <= '0';
                when 5924 => sda_i <= '0';
                when 5925 => sda_i <= '0';
                when 5926 => sda_i <= '0';
                when 5927 => sda_i <= '0';
                when 5928 => sda_i <= '0';
                when 5929 => sda_i <= '0';
                when 5930 => sda_i <= '0';
                when 5931 => sda_i <= '0';
                when 5932 => sda_i <= '0';
                when 5933 => sda_i <= '0';
                when 5934 => sda_i <= '0';
                when 5935 => sda_i <= '0';
                when 5936 => sda_i <= '0';
                when 5937 => sda_i <= '0';
                when 5938 => sda_i <= '1';
                when 5939 => sda_i <= '1';
                when 5940 => sda_i <= '0';
                when 5941 => sda_i <= '0';
                when 5942 => sda_i <= '0';
                when 5943 => sda_i <= '0';
                when 5944 => sda_i <= '0';
                when 5945 => sda_i <= '0';
                when 5946 => sda_i <= '0';
                when 5947 => sda_i <= '0';
                when 5948 => sda_i <= '0';
                when 5949 => sda_i <= '0';
                when 5950 => sda_i <= '0';
                when 5951 => sda_i <= '0';
                when 5952 => sda_i <= '0';
                when 5953 => sda_i <= '0';
                when 5954 => sda_i <= '0';
                when 5955 => sda_i <= '0';
                when 5956 => sda_i <= '0';
                when 5957 => sda_i <= '0';
                when 5958 => sda_i <= '0';
                when 5959 => sda_i <= '0';
                when 5960 => sda_i <= '0';
                when 5961 => sda_i <= '0';
                when 5962 => sda_i <= '0';
                when 5963 => sda_i <= '0';
                when 5964 => sda_i <= '0';
                when 5965 => sda_i <= '0';
                when 5966 => sda_i <= '0';
                when 5967 => sda_i <= '0';
                when 5968 => sda_i <= '0';
                when 5969 => sda_i <= '0';
                when 5970 => sda_i <= '0';
                when 5971 => sda_i <= '0';
                when 5972 => sda_i <= '0';
                when 5973 => sda_i <= '0';
                when 5974 => sda_i <= '0';
                when 5975 => sda_i <= '0';
                when 5976 => sda_i <= '0';
                when 5977 => sda_i <= '0';
                when 5978 => sda_i <= '0';
                when 5979 => sda_i <= '0';
                when 5980 => sda_i <= '0';
                when 5981 => sda_i <= '0';
                when 5982 => sda_i <= '0';
                when 5983 => sda_i <= '0';
                when 5984 => sda_i <= '0';
                when 5985 => sda_i <= '0';
                when 5986 => sda_i <= '0';
                when 5987 => sda_i <= '0';
                when 5988 => sda_i <= '0';
                when 5989 => sda_i <= '0';
                when 5990 => sda_i <= '0';
                when 5991 => sda_i <= '0';
                when 5992 => sda_i <= '0';
                when 5993 => sda_i <= '0';
                when 5994 => sda_i <= '0';
                when 5995 => sda_i <= '0';
                when 5996 => sda_i <= '0';
                when 5997 => sda_i <= '0';
                when 5998 => sda_i <= '0';
                when 5999 => sda_i <= '0';
                when 6000 => sda_i <= '0';
                when 6001 => sda_i <= '0';
                when 6002 => sda_i <= '0';
                when 6003 => sda_i <= '0';
                when 6004 => sda_i <= '0';
                when 6005 => sda_i <= '0';
                when 6006 => sda_i <= '0';
                when 6007 => sda_i <= '0';
                when 6008 => sda_i <= '0';
                when 6009 => sda_i <= '0';
                when 6010 => sda_i <= '0';
                when 6011 => sda_i <= '0';
                when 6012 => sda_i <= '0';
                when 6013 => sda_i <= '0';
                when 6014 => sda_i <= '0';
                when 6015 => sda_i <= '0';
                when 6016 => sda_i <= '0';
                when 6017 => sda_i <= '0';
                when 6018 => sda_i <= '0';
                when 6019 => sda_i <= '0';
                when 6020 => sda_i <= '0';
                when 6021 => sda_i <= '0';
                when 6022 => sda_i <= '0';
                when 6023 => sda_i <= '0';
                when 6024 => sda_i <= '0';
                when 6025 => sda_i <= '0';
                when 6026 => sda_i <= '0';
                when 6027 => sda_i <= '0';
                when 6028 => sda_i <= '0';
                when 6029 => sda_i <= '0';
                when 6030 => sda_i <= '0';
                when 6031 => sda_i <= '0';
                when 6032 => sda_i <= '0';
                when 6033 => sda_i <= '0';
                when 6034 => sda_i <= '0';
                when 6035 => sda_i <= '0';
                when 6036 => sda_i <= '0';
                when 6037 => sda_i <= '0';
                when 6038 => sda_i <= '0';
                when 6039 => sda_i <= '0';
                when 6040 => sda_i <= '0';
                when 6041 => sda_i <= '0';
                when 6042 => sda_i <= '0';
                when 6043 => sda_i <= '0';
                when 6044 => sda_i <= '0';
                when 6045 => sda_i <= '0';
                when 6046 => sda_i <= '1';
                when 6047 => sda_i <= '1';
                when 6048 => sda_i <= '0';
                when 6049 => sda_i <= '0';
                when 6050 => sda_i <= '0';
                when 6051 => sda_i <= '0';
                when 6052 => sda_i <= '0';
                when 6053 => sda_i <= '0';
                when 6054 => sda_i <= '0';
                when 6055 => sda_i <= '0';
                when 6056 => sda_i <= '0';
                when 6057 => sda_i <= '0';
                when 6058 => sda_i <= '0';
                when 6059 => sda_i <= '0';
                when 6060 => sda_i <= '0';
                when 6061 => sda_i <= '0';
                when 6062 => sda_i <= '0';
                when 6063 => sda_i <= '0';
                when 6064 => sda_i <= '0';
                when 6065 => sda_i <= '0';
                when 6066 => sda_i <= '0';
                when 6067 => sda_i <= '0';
                when 6068 => sda_i <= '0';
                when 6069 => sda_i <= '0';
                when 6070 => sda_i <= '0';
                when 6071 => sda_i <= '0';
                when 6072 => sda_i <= '0';
                when 6073 => sda_i <= '0';
                when 6074 => sda_i <= '0';
                when 6075 => sda_i <= '0';
                when 6076 => sda_i <= '0';
                when 6077 => sda_i <= '0';
                when 6078 => sda_i <= '0';
                when 6079 => sda_i <= '0';
                when 6080 => sda_i <= '0';
                when 6081 => sda_i <= '0';
                when 6082 => sda_i <= '0';
                when 6083 => sda_i <= '0';
                when 6084 => sda_i <= '0';
                when 6085 => sda_i <= '0';
                when 6086 => sda_i <= '0';
                when 6087 => sda_i <= '0';
                when 6088 => sda_i <= '0';
                when 6089 => sda_i <= '0';
                when 6090 => sda_i <= '0';
                when 6091 => sda_i <= '0';
                when 6092 => sda_i <= '0';
                when 6093 => sda_i <= '0';
                when 6094 => sda_i <= '0';
                when 6095 => sda_i <= '0';
                when 6096 => sda_i <= '0';
                when 6097 => sda_i <= '0';
                when 6098 => sda_i <= '0';
                when 6099 => sda_i <= '0';
                when 6100 => sda_i <= '0';
                when 6101 => sda_i <= '0';
                when 6102 => sda_i <= '0';
                when 6103 => sda_i <= '0';
                when 6104 => sda_i <= '0';
                when 6105 => sda_i <= '0';
                when 6106 => sda_i <= '0';
                when 6107 => sda_i <= '0';
                when 6108 => sda_i <= '0';
                when 6109 => sda_i <= '0';
                when 6110 => sda_i <= '0';
                when 6111 => sda_i <= '0';
                when 6112 => sda_i <= '0';
                when 6113 => sda_i <= '0';
                when 6114 => sda_i <= '0';
                when 6115 => sda_i <= '0';
                when 6116 => sda_i <= '0';
                when 6117 => sda_i <= '0';
                when 6118 => sda_i <= '0';
                when 6119 => sda_i <= '0';
                when 6120 => sda_i <= '0';
                when 6121 => sda_i <= '0';
                when 6122 => sda_i <= '0';
                when 6123 => sda_i <= '0';
                when 6124 => sda_i <= '0';
                when 6125 => sda_i <= '0';
                when 6126 => sda_i <= '0';
                when 6127 => sda_i <= '0';
                when 6128 => sda_i <= '0';
                when 6129 => sda_i <= '0';
                when 6130 => sda_i <= '0';
                when 6131 => sda_i <= '0';
                when 6132 => sda_i <= '0';
                when 6133 => sda_i <= '0';
                when 6134 => sda_i <= '0';
                when 6135 => sda_i <= '0';
                when 6136 => sda_i <= '0';
                when 6137 => sda_i <= '0';
                when 6138 => sda_i <= '0';
                when 6139 => sda_i <= '0';
                when 6140 => sda_i <= '0';
                when 6141 => sda_i <= '0';
                when 6142 => sda_i <= '0';
                when 6143 => sda_i <= '0';
                when 6144 => sda_i <= '0';
                when 6145 => sda_i <= '0';
                when 6146 => sda_i <= '0';
                when 6147 => sda_i <= '0';
                when 6148 => sda_i <= '0';
                when 6149 => sda_i <= '0';
                when 6150 => sda_i <= '0';
                when 6151 => sda_i <= '0';
                when 6152 => sda_i <= '0';
                when 6153 => sda_i <= '0';
                when 6154 => sda_i <= '1';
                when 6155 => sda_i <= '1';
                when 6156 => sda_i <= '0';
                when 6157 => sda_i <= '0';
                when 6158 => sda_i <= '0';
                when 6159 => sda_i <= '0';
                when 6160 => sda_i <= '0';
                when 6161 => sda_i <= '0';
                when 6162 => sda_i <= '0';
                when 6163 => sda_i <= '0';
                when 6164 => sda_i <= '0';
                when 6165 => sda_i <= '0';
                when 6166 => sda_i <= '0';
                when 6167 => sda_i <= '0';
                when 6168 => sda_i <= '0';
                when 6169 => sda_i <= '0';
                when 6170 => sda_i <= '0';
                when 6171 => sda_i <= '0';
                when 6172 => sda_i <= '0';
                when 6173 => sda_i <= '0';
                when 6174 => sda_i <= '0';
                when 6175 => sda_i <= '0';
                when 6176 => sda_i <= '0';
                when 6177 => sda_i <= '0';
                when 6178 => sda_i <= '0';
                when 6179 => sda_i <= '0';
                when 6180 => sda_i <= '0';
                when 6181 => sda_i <= '0';
                when 6182 => sda_i <= '0';
                when 6183 => sda_i <= '0';
                when 6184 => sda_i <= '0';
                when 6185 => sda_i <= '0';
                when 6186 => sda_i <= '0';
                when 6187 => sda_i <= '0';
                when 6188 => sda_i <= '0';
                when 6189 => sda_i <= '0';
                when 6190 => sda_i <= '0';
                when 6191 => sda_i <= '0';
                when 6192 => sda_i <= '0';
                when 6193 => sda_i <= '0';
                when 6194 => sda_i <= '0';
                when 6195 => sda_i <= '0';
                when 6196 => sda_i <= '0';
                when 6197 => sda_i <= '0';
                when 6198 => sda_i <= '0';
                when 6199 => sda_i <= '0';
                when 6200 => sda_i <= '0';
                when 6201 => sda_i <= '0';
                when 6202 => sda_i <= '0';
                when 6203 => sda_i <= '0';
                when 6204 => sda_i <= '0';
                when 6205 => sda_i <= '0';
                when 6206 => sda_i <= '0';
                when 6207 => sda_i <= '0';
                when 6208 => sda_i <= '0';
                when 6209 => sda_i <= '0';
                when 6210 => sda_i <= '0';
                when 6211 => sda_i <= '0';
                when 6212 => sda_i <= '0';
                when 6213 => sda_i <= '0';
                when 6214 => sda_i <= '0';
                when 6215 => sda_i <= '0';
                when 6216 => sda_i <= '0';
                when 6217 => sda_i <= '0';
                when 6218 => sda_i <= '0';
                when 6219 => sda_i <= '0';
                when 6220 => sda_i <= '0';
                when 6221 => sda_i <= '0';
                when 6222 => sda_i <= '0';
                when 6223 => sda_i <= '0';
                when 6224 => sda_i <= '0';
                when 6225 => sda_i <= '0';
                when 6226 => sda_i <= '0';
                when 6227 => sda_i <= '0';
                when 6228 => sda_i <= '0';
                when 6229 => sda_i <= '0';
                when 6230 => sda_i <= '0';
                when 6231 => sda_i <= '0';
                when 6232 => sda_i <= '0';
                when 6233 => sda_i <= '0';
                when 6234 => sda_i <= '0';
                when 6235 => sda_i <= '0';
                when 6236 => sda_i <= '0';
                when 6237 => sda_i <= '0';
                when 6238 => sda_i <= '0';
                when 6239 => sda_i <= '0';
                when 6240 => sda_i <= '0';
                when 6241 => sda_i <= '0';
                when 6242 => sda_i <= '0';
                when 6243 => sda_i <= '0';
                when 6244 => sda_i <= '0';
                when 6245 => sda_i <= '0';
                when 6246 => sda_i <= '0';
                when 6247 => sda_i <= '0';
                when 6248 => sda_i <= '0';
                when 6249 => sda_i <= '0';
                when 6250 => sda_i <= '0';
                when 6251 => sda_i <= '0';
                when 6252 => sda_i <= '0';
                when 6253 => sda_i <= '0';
                when 6254 => sda_i <= '0';
                when 6255 => sda_i <= '0';
                when 6256 => sda_i <= '0';
                when 6257 => sda_i <= '0';
                when 6258 => sda_i <= '0';
                when 6259 => sda_i <= '0';
                when 6260 => sda_i <= '0';
                when 6261 => sda_i <= '0';
                when 6262 => sda_i <= '1';
                when 6263 => sda_i <= '1';
                when 6264 => sda_i <= '0';
                when 6265 => sda_i <= '0';
                when 6266 => sda_i <= '0';
                when 6267 => sda_i <= '0';
                when 6268 => sda_i <= '0';
                when 6269 => sda_i <= '0';
                when 6270 => sda_i <= '0';
                when 6271 => sda_i <= '0';
                when 6272 => sda_i <= '0';
                when 6273 => sda_i <= '0';
                when 6274 => sda_i <= '0';
                when 6275 => sda_i <= '0';
                when 6276 => sda_i <= '0';
                when 6277 => sda_i <= '0';
                when 6278 => sda_i <= '0';
                when 6279 => sda_i <= '0';
                when 6280 => sda_i <= '0';
                when 6281 => sda_i <= '0';
                when 6282 => sda_i <= '0';
                when 6283 => sda_i <= '0';
                when 6284 => sda_i <= '0';
                when 6285 => sda_i <= '0';
                when 6286 => sda_i <= '0';
                when 6287 => sda_i <= '0';
                when 6288 => sda_i <= '0';
                when 6289 => sda_i <= '0';
                when 6290 => sda_i <= '0';
                when 6291 => sda_i <= '0';
                when 6292 => sda_i <= '0';
                when 6293 => sda_i <= '0';
                when 6294 => sda_i <= '0';
                when 6295 => sda_i <= '0';
                when 6296 => sda_i <= '0';
                when 6297 => sda_i <= '0';
                when 6298 => sda_i <= '0';
                when 6299 => sda_i <= '0';
                when 6300 => sda_i <= '0';
                when 6301 => sda_i <= '0';
                when 6302 => sda_i <= '0';
                when 6303 => sda_i <= '0';
                when 6304 => sda_i <= '0';
                when 6305 => sda_i <= '0';
                when 6306 => sda_i <= '0';
                when 6307 => sda_i <= '0';
                when 6308 => sda_i <= '0';
                when 6309 => sda_i <= '0';
                when 6310 => sda_i <= '0';
                when 6311 => sda_i <= '0';
                when 6312 => sda_i <= '0';
                when 6313 => sda_i <= '0';
                when 6314 => sda_i <= '0';
                when 6315 => sda_i <= '0';
                when 6316 => sda_i <= '0';
                when 6317 => sda_i <= '0';
                when 6318 => sda_i <= '0';
                when 6319 => sda_i <= '0';
                when 6320 => sda_i <= '0';
                when 6321 => sda_i <= '0';
                when 6322 => sda_i <= '0';
                when 6323 => sda_i <= '0';
                when 6324 => sda_i <= '0';
                when 6325 => sda_i <= '0';
                when 6326 => sda_i <= '0';
                when 6327 => sda_i <= '0';
                when 6328 => sda_i <= '0';
                when 6329 => sda_i <= '0';
                when 6330 => sda_i <= '0';
                when 6331 => sda_i <= '0';
                when 6332 => sda_i <= '0';
                when 6333 => sda_i <= '0';
                when 6334 => sda_i <= '0';
                when 6335 => sda_i <= '0';
                when 6336 => sda_i <= '0';
                when 6337 => sda_i <= '0';
                when 6338 => sda_i <= '0';
                when 6339 => sda_i <= '0';
                when 6340 => sda_i <= '0';
                when 6341 => sda_i <= '0';
                when 6342 => sda_i <= '0';
                when 6343 => sda_i <= '0';
                when 6344 => sda_i <= '0';
                when 6345 => sda_i <= '0';
                when 6346 => sda_i <= '0';
                when 6347 => sda_i <= '0';
                when 6348 => sda_i <= '0';
                when 6349 => sda_i <= '0';
                when 6350 => sda_i <= '0';
                when 6351 => sda_i <= '0';
                when 6352 => sda_i <= '0';
                when 6353 => sda_i <= '0';
                when 6354 => sda_i <= '0';
                when 6355 => sda_i <= '0';
                when 6356 => sda_i <= '0';
                when 6357 => sda_i <= '0';
                when 6358 => sda_i <= '0';
                when 6359 => sda_i <= '0';
                when 6360 => sda_i <= '0';
                when 6361 => sda_i <= '0';
                when 6362 => sda_i <= '0';
                when 6363 => sda_i <= '0';
                when 6364 => sda_i <= '0';
                when 6365 => sda_i <= '0';
                when 6366 => sda_i <= '0';
                when 6367 => sda_i <= '0';
                when 6368 => sda_i <= '0';
                when 6369 => sda_i <= '0';
                when 6370 => sda_i <= '1';
                when 6371 => sda_i <= '1';
                when 6372 => sda_i <= '1';
                when 6373 => sda_i <= '1';
                when 6374 => sda_i <= '1';
                when 6375 => sda_i <= '1';
                when 6376 => sda_i <= '1';
                when 6377 => sda_i <= '1';
                when 6378 => sda_i <= '1';
                when 6379 => sda_i <= '1';
                when 6380 => sda_i <= '1';
                when 6381 => sda_i <= '1';
                when 6382 => sda_i <= '1';
                when 6383 => sda_i <= '1';
                when 6384 => sda_i <= '0';
                when 6385 => sda_i <= '0';
                when 6386 => sda_i <= '0';
                when 6387 => sda_i <= '0';
                when 6388 => sda_i <= '0';
                when 6389 => sda_i <= '0';
                when 6390 => sda_i <= '0';
                when 6391 => sda_i <= '0';
                when 6392 => sda_i <= '0';
                when 6393 => sda_i <= '0';
                when 6394 => sda_i <= '0';
                when 6395 => sda_i <= '0';
                when 6396 => sda_i <= '1';
                when 6397 => sda_i <= '1';
                when 6398 => sda_i <= '1';
                when 6399 => sda_i <= '1';
                when 6400 => sda_i <= '1';
                when 6401 => sda_i <= '1';
                when 6402 => sda_i <= '1';
                when 6403 => sda_i <= '1';
                when 6404 => sda_i <= '1';
                when 6405 => sda_i <= '1';
                when 6406 => sda_i <= '1';
                when 6407 => sda_i <= '1';
                when 6408 => sda_i <= '1';
                when 6409 => sda_i <= '1';
                when 6410 => sda_i <= '1';
                when 6411 => sda_i <= '1';
                when 6412 => sda_i <= '1';
                when 6413 => sda_i <= '1';
                when 6414 => sda_i <= '1';
                when 6415 => sda_i <= '1';
                when 6416 => sda_i <= '1';
                when 6417 => sda_i <= '1';
                when 6418 => sda_i <= '1';
                when 6419 => sda_i <= '1';
                when 6420 => sda_i <= '1';
                when 6421 => sda_i <= '1';
                when 6422 => sda_i <= '1';
                when 6423 => sda_i <= '1';
                when 6424 => sda_i <= '1';
                when 6425 => sda_i <= '1';
                when 6426 => sda_i <= '1';
                when 6427 => sda_i <= '1';
                when 6428 => sda_i <= '1';
                when 6429 => sda_i <= '1';
                when 6430 => sda_i <= '1';
                when 6431 => sda_i <= '1';
                when 6432 => sda_i <= '1';
                when 6433 => sda_i <= '1';
                when 6434 => sda_i <= '1';
                when 6435 => sda_i <= '1';
                when 6436 => sda_i <= '1';
                when 6437 => sda_i <= '1';
                when 6438 => sda_i <= '1';
                when 6439 => sda_i <= '1';
                when 6440 => sda_i <= '1';
                when 6441 => sda_i <= '1';
                when 6442 => sda_i <= '1';
                when 6443 => sda_i <= '1';
                when 6444 => sda_i <= '1';
                when 6445 => sda_i <= '1';
                when 6446 => sda_i <= '1';
                when 6447 => sda_i <= '1';
                when 6448 => sda_i <= '1';
                when 6449 => sda_i <= '1';
                when 6450 => sda_i <= '1';
                when 6451 => sda_i <= '1';
                when 6452 => sda_i <= '1';
                when 6453 => sda_i <= '1';
                when 6454 => sda_i <= '1';
                when 6455 => sda_i <= '1';
                when 6456 => sda_i <= '1';
                when 6457 => sda_i <= '1';
                when 6458 => sda_i <= '1';
                when 6459 => sda_i <= '1';
                when 6460 => sda_i <= '1';
                when 6461 => sda_i <= '1';
                when 6462 => sda_i <= '1';
                when 6463 => sda_i <= '1';
                when 6464 => sda_i <= '1';
                when 6465 => sda_i <= '1';
                when 6466 => sda_i <= '1';
                when 6467 => sda_i <= '1';
                when 6468 => sda_i <= '1';
                when 6469 => sda_i <= '1';
                when 6470 => sda_i <= '1';
                when 6471 => sda_i <= '1';
                when 6472 => sda_i <= '1';
                when 6473 => sda_i <= '1';
                when 6474 => sda_i <= '1';
                when 6475 => sda_i <= '1';
                when 6476 => sda_i <= '1';
                when 6477 => sda_i <= '1';
                when 6478 => sda_i <= '1';
                when 6479 => sda_i <= '1';
                when 6480 => sda_i <= '1';
                when 6481 => sda_i <= '1';
                when 6482 => sda_i <= '1';
                when 6483 => sda_i <= '1';
                when 6484 => sda_i <= '1';
                when 6485 => sda_i <= '1';
                when 6486 => sda_i <= '1';
                when 6487 => sda_i <= '1';
                when 6488 => sda_i <= '1';
                when 6489 => sda_i <= '1';
                when 6490 => sda_i <= '1';
                when 6491 => sda_i <= '1';
                when 6492 => sda_i <= '1';
                when 6493 => sda_i <= '1';
                when 6494 => sda_i <= '1';
                when 6495 => sda_i <= '1';
                when 6496 => sda_i <= '1';
                when 6497 => sda_i <= '1';
                when 6498 => sda_i <= '1';
                when 6499 => sda_i <= '1';
                when 6500 => sda_i <= '1';
                when 6501 => sda_i <= '1';
                when 6502 => sda_i <= '1';
                when 6503 => sda_i <= '1';
                when 6504 => sda_i <= '1';
                when 6505 => sda_i <= '1';
                when 6506 => sda_i <= '1';
                when 6507 => sda_i <= '1';
                when 6508 => sda_i <= '1';
                when 6509 => sda_i <= '1';
                when 6510 => sda_i <= '1';
                when 6511 => sda_i <= '1';
                when 6512 => sda_i <= '1';
                when 6513 => sda_i <= '1';
                when 6514 => sda_i <= '1';
                when 6515 => sda_i <= '1';
                when 6516 => sda_i <= '1';
                when 6517 => sda_i <= '1';
                when 6518 => sda_i <= '1';
                when 6519 => sda_i <= '1';
                when 6520 => sda_i <= '1';
                when 6521 => sda_i <= '1';
                when 6522 => sda_i <= '1';
                when 6523 => sda_i <= '1';
                when 6524 => sda_i <= '1';
                when 6525 => sda_i <= '1';
                when 6526 => sda_i <= '1';
                when 6527 => sda_i <= '1';
                when 6528 => sda_i <= '1';
                when 6529 => sda_i <= '1';
                when 6530 => sda_i <= '1';
                when 6531 => sda_i <= '1';
                when 6532 => sda_i <= '1';
                when 6533 => sda_i <= '1';
                when 6534 => sda_i <= '1';
                when 6535 => sda_i <= '1';
                when 6536 => sda_i <= '1';
                when 6537 => sda_i <= '1';
                when 6538 => sda_i <= '1';
                when 6539 => sda_i <= '1';
                when 6540 => sda_i <= '1';
                when 6541 => sda_i <= '1';
                when 6542 => sda_i <= '1';
                when 6543 => sda_i <= '1';
                when 6544 => sda_i <= '1';
                when 6545 => sda_i <= '1';
                when 6546 => sda_i <= '1';
                when 6547 => sda_i <= '1';
                when 6548 => sda_i <= '1';
                when 6549 => sda_i <= '1';
                when 6550 => sda_i <= '1';
                when 6551 => sda_i <= '1';
                when 6552 => sda_i <= '1';
                when 6553 => sda_i <= '1';
                when 6554 => sda_i <= '1';
                when 6555 => sda_i <= '1';
                when 6556 => sda_i <= '1';
                when 6557 => sda_i <= '1';
                when 6558 => sda_i <= '1';
                when 6559 => sda_i <= '1';
                when 6560 => sda_i <= '1';
                when 6561 => sda_i <= '1';
                when 6562 => sda_i <= '1';
                when 6563 => sda_i <= '1';
                when 6564 => sda_i <= '1';
                when 6565 => sda_i <= '1';
                when 6566 => sda_i <= '1';
                when 6567 => sda_i <= '1';
                when 6568 => sda_i <= '1';
                when 6569 => sda_i <= '1';
                when 6570 => sda_i <= '1';
                when 6571 => sda_i <= '1';
                when 6572 => sda_i <= '1';
                when 6573 => sda_i <= '1';
                when 6574 => sda_i <= '1';
                when 6575 => sda_i <= '1';
                when 6576 => sda_i <= '1';
                when 6577 => sda_i <= '1';
                when 6578 => sda_i <= '1';
                when 6579 => sda_i <= '1';
                when 6580 => sda_i <= '1';
                when 6581 => sda_i <= '1';
                when 6582 => sda_i <= '1';
                when 6583 => sda_i <= '1';
                when 6584 => sda_i <= '1';
                when 6585 => sda_i <= '1';
                when 6586 => sda_i <= '1';
                when 6587 => sda_i <= '1';
                when 6588 => sda_i <= '1';
                when 6589 => sda_i <= '1';
                when 6590 => sda_i <= '1';
                when 6591 => sda_i <= '1';
                when 6592 => sda_i <= '1';
                when 6593 => sda_i <= '1';
                when 6594 => sda_i <= '1';
                when 6595 => sda_i <= '1';
                when 6596 => sda_i <= '1';
                when 6597 => sda_i <= '1';
                when 6598 => sda_i <= '1';
                when 6599 => sda_i <= '1';
                when 6600 => sda_i <= '1';
                when 6601 => sda_i <= '1';
                when 6602 => sda_i <= '1';
                when 6603 => sda_i <= '1';
                when 6604 => sda_i <= '1';
                when 6605 => sda_i <= '1';
                when 6606 => sda_i <= '1';
                when 6607 => sda_i <= '1';
                when 6608 => sda_i <= '1';
                when 6609 => sda_i <= '1';
                when 6610 => sda_i <= '1';
                when 6611 => sda_i <= '1';
                when 6612 => sda_i <= '1';
                when 6613 => sda_i <= '1';
                when 6614 => sda_i <= '1';
                when 6615 => sda_i <= '1';
                when 6616 => sda_i <= '1';
                when 6617 => sda_i <= '1';
                when 6618 => sda_i <= '1';
                when 6619 => sda_i <= '1';
                when 6620 => sda_i <= '1';
                when 6621 => sda_i <= '1';
                when 6622 => sda_i <= '1';
                when 6623 => sda_i <= '1';
                when 6624 => sda_i <= '1';
                when 6625 => sda_i <= '1';
                when 6626 => sda_i <= '1';
                when 6627 => sda_i <= '1';
                when 6628 => sda_i <= '1';
                when 6629 => sda_i <= '1';
                when 6630 => sda_i <= '1';
                when 6631 => sda_i <= '1';
                when 6632 => sda_i <= '1';
                when 6633 => sda_i <= '1';
                when 6634 => sda_i <= '1';
                when 6635 => sda_i <= '1';
                when 6636 => sda_i <= '1';
                when 6637 => sda_i <= '1';
                when 6638 => sda_i <= '1';
                when 6639 => sda_i <= '1';
                when 6640 => sda_i <= '1';
                when 6641 => sda_i <= '1';
                when 6642 => sda_i <= '1';
                when 6643 => sda_i <= '1';
                when 6644 => sda_i <= '1';
                when 6645 => sda_i <= '1';
                when 6646 => sda_i <= '1';
                when 6647 => sda_i <= '1';
                when 6648 => sda_i <= '1';
                when 6649 => sda_i <= '1';
                when 6650 => sda_i <= '1';
                when 6651 => sda_i <= '1';
                when 6652 => sda_i <= '1';
                when 6653 => sda_i <= '1';
                when 6654 => sda_i <= '1';
                when 6655 => sda_i <= '1';
                when 6656 => sda_i <= '1';
                when 6657 => sda_i <= '1';
                when 6658 => sda_i <= '1';
                when 6659 => sda_i <= '1';
                when 6660 => sda_i <= '1';
                when 6661 => sda_i <= '1';
                when 6662 => sda_i <= '1';
                when 6663 => sda_i <= '1';
                when 6664 => sda_i <= '1';
                when 6665 => sda_i <= '1';
                when 6666 => sda_i <= '1';
                when 6667 => sda_i <= '1';
                when 6668 => sda_i <= '1';
                when 6669 => sda_i <= '1';
                when 6670 => sda_i <= '1';
                when 6671 => sda_i <= '1';
                when 6672 => sda_i <= '1';
                when 6673 => sda_i <= '1';
                when 6674 => sda_i <= '1';
                when 6675 => sda_i <= '1';
                when 6676 => sda_i <= '1';
                when 6677 => sda_i <= '1';
                when 6678 => sda_i <= '1';
                when 6679 => sda_i <= '1';
                when 6680 => sda_i <= '1';
                when 6681 => sda_i <= '1';
                when 6682 => sda_i <= '1';
                when 6683 => sda_i <= '1';
                when 6684 => sda_i <= '1';
                when 6685 => sda_i <= '1';
                when 6686 => sda_i <= '1';
                when 6687 => sda_i <= '1';
                when 6688 => sda_i <= '1';
                when 6689 => sda_i <= '1';
                when 6690 => sda_i <= '1';
                when 6691 => sda_i <= '1';
                when 6692 => sda_i <= '1';
                when 6693 => sda_i <= '1';
                when 6694 => sda_i <= '1';
                when 6695 => sda_i <= '1';
                when 6696 => sda_i <= '1';
                when 6697 => sda_i <= '1';
                when 6698 => sda_i <= '1';
                when 6699 => sda_i <= '1';
                when 6700 => sda_i <= '1';
                when 6701 => sda_i <= '1';
                when 6702 => sda_i <= '1';
                when 6703 => sda_i <= '1';
                when 6704 => sda_i <= '1';
                when 6705 => sda_i <= '1';
                when 6706 => sda_i <= '1';
                when 6707 => sda_i <= '1';
                when 6708 => sda_i <= '1';
                when 6709 => sda_i <= '1';
                when 6710 => sda_i <= '1';
                when 6711 => sda_i <= '1';
                when 6712 => sda_i <= '1';
                when 6713 => sda_i <= '1';
                when 6714 => sda_i <= '1';
                when 6715 => sda_i <= '1';
                when 6716 => sda_i <= '1';
                when 6717 => sda_i <= '1';
                when 6718 => sda_i <= '1';
                when 6719 => sda_i <= '1';
                when 6720 => sda_i <= '1';
                when 6721 => sda_i <= '1';
                when 6722 => sda_i <= '1';
                when 6723 => sda_i <= '1';
                when 6724 => sda_i <= '1';
                when 6725 => sda_i <= '1';
                when 6726 => sda_i <= '1';
                when 6727 => sda_i <= '1';
                when 6728 => sda_i <= '1';
                when 6729 => sda_i <= '1';
                when 6730 => sda_i <= '1';
                when 6731 => sda_i <= '1';
                when 6732 => sda_i <= '1';
                when 6733 => sda_i <= '1';
                when 6734 => sda_i <= '1';
                when 6735 => sda_i <= '1';
                when 6736 => sda_i <= '1';
                when 6737 => sda_i <= '1';
                when 6738 => sda_i <= '1';
                when 6739 => sda_i <= '1';
                when 6740 => sda_i <= '1';
                when 6741 => sda_i <= '1';
                when 6742 => sda_i <= '1';
                when 6743 => sda_i <= '1';
                when 6744 => sda_i <= '1';
                when 6745 => sda_i <= '1';
                when 6746 => sda_i <= '1';
                when 6747 => sda_i <= '1';
                when 6748 => sda_i <= '1';
                when 6749 => sda_i <= '1';
                when 6750 => sda_i <= '1';
                when 6751 => sda_i <= '1';
                when 6752 => sda_i <= '1';
                when 6753 => sda_i <= '1';
                when 6754 => sda_i <= '1';
                when 6755 => sda_i <= '1';
                when 6756 => sda_i <= '1';
                when 6757 => sda_i <= '1';
                when 6758 => sda_i <= '1';
                when 6759 => sda_i <= '1';
                when 6760 => sda_i <= '1';
                when 6761 => sda_i <= '1';
                when 6762 => sda_i <= '1';
                when 6763 => sda_i <= '1';
                when 6764 => sda_i <= '1';
                when 6765 => sda_i <= '1';
                when 6766 => sda_i <= '1';
                when 6767 => sda_i <= '1';
                when 6768 => sda_i <= '1';
                when 6769 => sda_i <= '1';
                when 6770 => sda_i <= '1';
                when 6771 => sda_i <= '1';
                when 6772 => sda_i <= '1';
                when 6773 => sda_i <= '1';
                when 6774 => sda_i <= '1';
                when 6775 => sda_i <= '1';
                when 6776 => sda_i <= '1';
                when 6777 => sda_i <= '1';
                when 6778 => sda_i <= '1';
                when 6779 => sda_i <= '1';
                when 6780 => sda_i <= '1';
                when 6781 => sda_i <= '1';
                when 6782 => sda_i <= '1';
                when 6783 => sda_i <= '1';
                when 6784 => sda_i <= '1';
                when 6785 => sda_i <= '1';
                when 6786 => sda_i <= '1';
                when 6787 => sda_i <= '1';
                when 6788 => sda_i <= '1';
                when 6789 => sda_i <= '1';
                when 6790 => sda_i <= '1';
                when 6791 => sda_i <= '1';
                when 6792 => sda_i <= '1';
                when 6793 => sda_i <= '1';
                when 6794 => sda_i <= '1';
                when 6795 => sda_i <= '1';
                when 6796 => sda_i <= '1';
                when 6797 => sda_i <= '1';
                when 6798 => sda_i <= '1';
                when 6799 => sda_i <= '1';
                when 6800 => sda_i <= '1';
                when 6801 => sda_i <= '1';
                when 6802 => sda_i <= '1';
                when 6803 => sda_i <= '1';
                when 6804 => sda_i <= '1';
                when 6805 => sda_i <= '1';
                when 6806 => sda_i <= '1';
                when 6807 => sda_i <= '1';
                when 6808 => sda_i <= '1';
                when 6809 => sda_i <= '1';
                when 6810 => sda_i <= '1';
                when 6811 => sda_i <= '1';
                when 6812 => sda_i <= '1';
                when 6813 => sda_i <= '1';
                when 6814 => sda_i <= '1';
                when 6815 => sda_i <= '1';
                when 6816 => sda_i <= '1';
                when 6817 => sda_i <= '1';
                when 6818 => sda_i <= '1';
                when 6819 => sda_i <= '1';
                when 6820 => sda_i <= '1';
                when 6821 => sda_i <= '1';
                when 6822 => sda_i <= '1';
                when 6823 => sda_i <= '1';
                when 6824 => sda_i <= '1';
                when 6825 => sda_i <= '1';
                when 6826 => sda_i <= '1';
                when 6827 => sda_i <= '1';
                when 6828 => sda_i <= '1';
                when 6829 => sda_i <= '1';
                when 6830 => sda_i <= '1';
                when 6831 => sda_i <= '1';
                when 6832 => sda_i <= '1';
                when 6833 => sda_i <= '1';
                when 6834 => sda_i <= '1';
                when 6835 => sda_i <= '1';
                when 6836 => sda_i <= '1';
                when 6837 => sda_i <= '1';
                when 6838 => sda_i <= '1';
                when 6839 => sda_i <= '1';
                when 6840 => sda_i <= '1';
                when 6841 => sda_i <= '1';
                when 6842 => sda_i <= '1';
                when 6843 => sda_i <= '1';
                when 6844 => sda_i <= '1';
                when 6845 => sda_i <= '1';
                when 6846 => sda_i <= '1';
                when 6847 => sda_i <= '1';
                when 6848 => sda_i <= '1';
                when 6849 => sda_i <= '1';
                when 6850 => sda_i <= '1';
                when 6851 => sda_i <= '1';
                when 6852 => sda_i <= '1';
                when 6853 => sda_i <= '1';
                when 6854 => sda_i <= '1';
                when 6855 => sda_i <= '1';
                when 6856 => sda_i <= '1';
                when 6857 => sda_i <= '1';
                when 6858 => sda_i <= '1';
                when 6859 => sda_i <= '1';
                when 6860 => sda_i <= '1';
                when 6861 => sda_i <= '1';
                when 6862 => sda_i <= '1';
                when 6863 => sda_i <= '1';
                when 6864 => sda_i <= '1';
                when 6865 => sda_i <= '1';
                when 6866 => sda_i <= '1';
                when 6867 => sda_i <= '1';
                when 6868 => sda_i <= '1';
                when 6869 => sda_i <= '1';
                when 6870 => sda_i <= '1';
                when 6871 => sda_i <= '1';
                when 6872 => sda_i <= '1';
                when 6873 => sda_i <= '1';
                when 6874 => sda_i <= '1';
                when 6875 => sda_i <= '1';
                when 6876 => sda_i <= '1';
                when 6877 => sda_i <= '1';
                when 6878 => sda_i <= '1';
                when 6879 => sda_i <= '1';
                when 6880 => sda_i <= '1';
                when 6881 => sda_i <= '1';
                when 6882 => sda_i <= '1';
                when 6883 => sda_i <= '1';
                when 6884 => sda_i <= '1';
                when 6885 => sda_i <= '1';
                when 6886 => sda_i <= '1';
                when 6887 => sda_i <= '1';
                when 6888 => sda_i <= '1';
                when 6889 => sda_i <= '1';
                when 6890 => sda_i <= '1';
                when 6891 => sda_i <= '1';
                when 6892 => sda_i <= '1';
                when 6893 => sda_i <= '1';
                when 6894 => sda_i <= '1';
                when 6895 => sda_i <= '1';
                when 6896 => sda_i <= '1';
                when 6897 => sda_i <= '1';
                when 6898 => sda_i <= '1';
                when 6899 => sda_i <= '1';
                when 6900 => sda_i <= '1';
                when 6901 => sda_i <= '1';
                when 6902 => sda_i <= '1';
                when 6903 => sda_i <= '1';
                when 6904 => sda_i <= '1';
                when 6905 => sda_i <= '1';
                when 6906 => sda_i <= '1';
                when 6907 => sda_i <= '1';
                when 6908 => sda_i <= '1';
                when 6909 => sda_i <= '1';
                when 6910 => sda_i <= '1';
                when 6911 => sda_i <= '1';
                when 6912 => sda_i <= '1';
                when 6913 => sda_i <= '1';
                when 6914 => sda_i <= '1';
                when 6915 => sda_i <= '1';
                when 6916 => sda_i <= '1';
                when 6917 => sda_i <= '1';
                when 6918 => sda_i <= '1';
                when 6919 => sda_i <= '1';
                when 6920 => sda_i <= '1';
                when 6921 => sda_i <= '1';
                when 6922 => sda_i <= '1';
                when 6923 => sda_i <= '1';
                when 6924 => sda_i <= '1';
                when 6925 => sda_i <= '1';
                when 6926 => sda_i <= '1';
                when 6927 => sda_i <= '1';
                when 6928 => sda_i <= '1';
                when 6929 => sda_i <= '1';
                when 6930 => sda_i <= '1';
                when 6931 => sda_i <= '1';
                when 6932 => sda_i <= '1';
                when 6933 => sda_i <= '1';
                when 6934 => sda_i <= '1';
                when 6935 => sda_i <= '1';
                when 6936 => sda_i <= '1';
                when 6937 => sda_i <= '1';
                when 6938 => sda_i <= '1';
                when 6939 => sda_i <= '1';
                when 6940 => sda_i <= '1';
                when 6941 => sda_i <= '1';
                when 6942 => sda_i <= '1';
                when 6943 => sda_i <= '1';
                when 6944 => sda_i <= '1';
                when 6945 => sda_i <= '1';
                when 6946 => sda_i <= '1';
                when 6947 => sda_i <= '1';
                when 6948 => sda_i <= '1';
                when 6949 => sda_i <= '1';
                when 6950 => sda_i <= '1';
                when 6951 => sda_i <= '1';
                when 6952 => sda_i <= '1';
                when 6953 => sda_i <= '1';
                when 6954 => sda_i <= '1';
                when 6955 => sda_i <= '1';
                when 6956 => sda_i <= '1';
                when 6957 => sda_i <= '1';
                when 6958 => sda_i <= '1';
                when 6959 => sda_i <= '1';
                when 6960 => sda_i <= '1';
                when 6961 => sda_i <= '1';
                when 6962 => sda_i <= '1';
                when 6963 => sda_i <= '1';
                when 6964 => sda_i <= '1';
                when 6965 => sda_i <= '1';
                when 6966 => sda_i <= '1';
                when 6967 => sda_i <= '1';
                when 6968 => sda_i <= '1';
                when 6969 => sda_i <= '1';
                when 6970 => sda_i <= '1';
                when 6971 => sda_i <= '1';
                when 6972 => sda_i <= '1';
                when 6973 => sda_i <= '1';
                when 6974 => sda_i <= '1';
                when 6975 => sda_i <= '1';
                when 6976 => sda_i <= '1';
                when 6977 => sda_i <= '1';
                when 6978 => sda_i <= '1';
                when 6979 => sda_i <= '1';
                when 6980 => sda_i <= '1';
                when 6981 => sda_i <= '1';
                when 6982 => sda_i <= '1';
                when 6983 => sda_i <= '1';
                when 6984 => sda_i <= '1';
                when 6985 => sda_i <= '1';
                when 6986 => sda_i <= '1';
                when 6987 => sda_i <= '1';
                when 6988 => sda_i <= '1';
                when 6989 => sda_i <= '1';
                when 6990 => sda_i <= '1';
                when 6991 => sda_i <= '1';
                when 6992 => sda_i <= '1';
                when 6993 => sda_i <= '1';
                when 6994 => sda_i <= '1';
                when 6995 => sda_i <= '1';
                when 6996 => sda_i <= '1';
                when 6997 => sda_i <= '1';
                when 6998 => sda_i <= '1';
                when 6999 => sda_i <= '1';
                when 7000 => sda_i <= '1';
                when 7001 => sda_i <= '1';
                when 7002 => sda_i <= '1';
                when 7003 => sda_i <= '1';
                when 7004 => sda_i <= '1';
                when 7005 => sda_i <= '1';
                when 7006 => sda_i <= '1';
                when 7007 => sda_i <= '1';
                when 7008 => sda_i <= '1';
                when 7009 => sda_i <= '1';
                when 7010 => sda_i <= '1';
                when 7011 => sda_i <= '1';
                when 7012 => sda_i <= '1';
                when 7013 => sda_i <= '1';
                when 7014 => sda_i <= '1';
                when 7015 => sda_i <= '1';
                when 7016 => sda_i <= '1';
                when 7017 => sda_i <= '1';
                when 7018 => sda_i <= '1';
                when 7019 => sda_i <= '1';
                when 7020 => sda_i <= '1';
                when 7021 => sda_i <= '1';
                when 7022 => sda_i <= '1';
                when 7023 => sda_i <= '1';
                when 7024 => sda_i <= '1';
                when 7025 => sda_i <= '1';
                when 7026 => sda_i <= '1';
                when 7027 => sda_i <= '1';
                when 7028 => sda_i <= '1';
                when 7029 => sda_i <= '1';
                when 7030 => sda_i <= '1';
                when 7031 => sda_i <= '1';
                when 7032 => sda_i <= '1';
                when 7033 => sda_i <= '1';
                when 7034 => sda_i <= '1';
                when 7035 => sda_i <= '1';
                when 7036 => sda_i <= '1';
                when 7037 => sda_i <= '1';
                when 7038 => sda_i <= '1';
                when 7039 => sda_i <= '1';
                when 7040 => sda_i <= '1';
                when 7041 => sda_i <= '1';
                when 7042 => sda_i <= '1';
                when 7043 => sda_i <= '1';
                when 7044 => sda_i <= '1';
                when 7045 => sda_i <= '1';
                when 7046 => sda_i <= '1';
                when 7047 => sda_i <= '1';
                when 7048 => sda_i <= '1';
                when 7049 => sda_i <= '1';
                when 7050 => sda_i <= '1';
                when 7051 => sda_i <= '1';
                when 7052 => sda_i <= '1';
                when 7053 => sda_i <= '1';
                when 7054 => sda_i <= '1';
                when 7055 => sda_i <= '1';
                when 7056 => sda_i <= '1';
                when 7057 => sda_i <= '1';
                when 7058 => sda_i <= '1';
                when 7059 => sda_i <= '1';
                when 7060 => sda_i <= '1';
                when 7061 => sda_i <= '1';
                when 7062 => sda_i <= '1';
                when 7063 => sda_i <= '1';
                when 7064 => sda_i <= '1';
                when 7065 => sda_i <= '1';
                when 7066 => sda_i <= '1';
                when 7067 => sda_i <= '1';
                when 7068 => sda_i <= '1';
                when 7069 => sda_i <= '1';
                when 7070 => sda_i <= '1';
                when 7071 => sda_i <= '1';
                when 7072 => sda_i <= '1';
                when 7073 => sda_i <= '1';
                when 7074 => sda_i <= '1';
                when 7075 => sda_i <= '1';
                when 7076 => sda_i <= '1';
                when 7077 => sda_i <= '1';
                when 7078 => sda_i <= '1';
                when 7079 => sda_i <= '1';
                when 7080 => sda_i <= '1';
                when 7081 => sda_i <= '1';
                when 7082 => sda_i <= '1';
                when 7083 => sda_i <= '1';
                when 7084 => sda_i <= '1';
                when 7085 => sda_i <= '1';
                when 7086 => sda_i <= '1';
                when 7087 => sda_i <= '1';
                when 7088 => sda_i <= '1';
                when 7089 => sda_i <= '1';
                when 7090 => sda_i <= '1';
                when 7091 => sda_i <= '1';
                when 7092 => sda_i <= '1';
                when 7093 => sda_i <= '1';
                when 7094 => sda_i <= '1';
                when 7095 => sda_i <= '1';
                when 7096 => sda_i <= '1';
                when 7097 => sda_i <= '1';
                when 7098 => sda_i <= '1';
                when 7099 => sda_i <= '1';
                when 7100 => sda_i <= '1';
                when 7101 => sda_i <= '1';
                when 7102 => sda_i <= '1';
                when 7103 => sda_i <= '1';
                when 7104 => sda_i <= '1';
                when 7105 => sda_i <= '1';
                when 7106 => sda_i <= '1';
                when 7107 => sda_i <= '1';
                when 7108 => sda_i <= '1';
                when 7109 => sda_i <= '1';
                when 7110 => sda_i <= '1';
                when 7111 => sda_i <= '1';
                when 7112 => sda_i <= '1';
                when 7113 => sda_i <= '1';
                when 7114 => sda_i <= '1';
                when 7115 => sda_i <= '1';
                when 7116 => sda_i <= '1';
                when 7117 => sda_i <= '1';
                when 7118 => sda_i <= '1';
                when 7119 => sda_i <= '1';
                when 7120 => sda_i <= '1';
                when 7121 => sda_i <= '1';
                when 7122 => sda_i <= '1';
                when 7123 => sda_i <= '1';
                when 7124 => sda_i <= '1';
                when 7125 => sda_i <= '1';
                when 7126 => sda_i <= '1';
                when 7127 => sda_i <= '1';
                when 7128 => sda_i <= '1';
                when 7129 => sda_i <= '1';
                when 7130 => sda_i <= '1';
                when 7131 => sda_i <= '1';
                when 7132 => sda_i <= '1';
                when 7133 => sda_i <= '1';
                when 7134 => sda_i <= '1';
                when 7135 => sda_i <= '1';
                when 7136 => sda_i <= '1';
                when 7137 => sda_i <= '1';
                when 7138 => sda_i <= '1';
                when 7139 => sda_i <= '1';
                when 7140 => sda_i <= '1';
                when 7141 => sda_i <= '1';
                when 7142 => sda_i <= '1';
                when 7143 => sda_i <= '1';
                when 7144 => sda_i <= '1';
                when 7145 => sda_i <= '1';
                when 7146 => sda_i <= '1';
                when 7147 => sda_i <= '1';
                when 7148 => sda_i <= '1';
                when 7149 => sda_i <= '1';
                when 7150 => sda_i <= '1';
                when 7151 => sda_i <= '1';
                when 7152 => sda_i <= '1';
                when 7153 => sda_i <= '1';
                when 7154 => sda_i <= '1';
                when 7155 => sda_i <= '1';
                when 7156 => sda_i <= '1';
                when 7157 => sda_i <= '1';
                when 7158 => sda_i <= '1';
                when 7159 => sda_i <= '1';
                when 7160 => sda_i <= '1';
                when 7161 => sda_i <= '1';
                when 7162 => sda_i <= '1';
                when 7163 => sda_i <= '1';
                when 7164 => sda_i <= '1';
                when 7165 => sda_i <= '1';
                when 7166 => sda_i <= '1';
                when 7167 => sda_i <= '1';
                when 7168 => sda_i <= '1';
                when 7169 => sda_i <= '1';
                when 7170 => sda_i <= '1';
                when 7171 => sda_i <= '1';
                when 7172 => sda_i <= '1';
                when 7173 => sda_i <= '1';
                when 7174 => sda_i <= '1';
                when 7175 => sda_i <= '1';
                when 7176 => sda_i <= '1';
                when 7177 => sda_i <= '1';
                when 7178 => sda_i <= '1';
                when 7179 => sda_i <= '1';
                when 7180 => sda_i <= '1';
                when 7181 => sda_i <= '1';
                when 7182 => sda_i <= '1';
                when 7183 => sda_i <= '1';
                when 7184 => sda_i <= '1';
                when 7185 => sda_i <= '1';
                when 7186 => sda_i <= '1';
                when 7187 => sda_i <= '1';
                when 7188 => sda_i <= '1';
                when 7189 => sda_i <= '1';
                when 7190 => sda_i <= '1';
                when 7191 => sda_i <= '1';
                when 7192 => sda_i <= '1';
                when 7193 => sda_i <= '1';
                when 7194 => sda_i <= '1';
                when 7195 => sda_i <= '1';
                when 7196 => sda_i <= '1';
                when 7197 => sda_i <= '1';
                when 7198 => sda_i <= '1';
                when 7199 => sda_i <= '1';
                when 7200 => sda_i <= '1';
                when 7201 => sda_i <= '1';
                when 7202 => sda_i <= '1';
                when 7203 => sda_i <= '1';
                when 7204 => sda_i <= '1';
                when 7205 => sda_i <= '1';
                when 7206 => sda_i <= '1';
                when 7207 => sda_i <= '1';
                when 7208 => sda_i <= '1';
                when 7209 => sda_i <= '1';
                when 7210 => sda_i <= '1';
                when 7211 => sda_i <= '1';
                when 7212 => sda_i <= '1';
                when 7213 => sda_i <= '1';
                when 7214 => sda_i <= '1';
                when 7215 => sda_i <= '1';
                when 7216 => sda_i <= '1';
                when 7217 => sda_i <= '1';
                when 7218 => sda_i <= '1';
                when 7219 => sda_i <= '1';
                when 7220 => sda_i <= '1';
                when 7221 => sda_i <= '1';
                when 7222 => sda_i <= '1';
                when 7223 => sda_i <= '1';
                when 7224 => sda_i <= '1';
                when 7225 => sda_i <= '1';
                when 7226 => sda_i <= '1';
                when 7227 => sda_i <= '1';
                when 7228 => sda_i <= '1';
                when 7229 => sda_i <= '1';
                when 7230 => sda_i <= '1';
                when 7231 => sda_i <= '1';
                when 7232 => sda_i <= '1';
                when 7233 => sda_i <= '1';
                when 7234 => sda_i <= '1';
                when 7235 => sda_i <= '1';
                when 7236 => sda_i <= '1';
                when 7237 => sda_i <= '1';
                when 7238 => sda_i <= '1';
                when 7239 => sda_i <= '1';
                when 7240 => sda_i <= '1';
                when 7241 => sda_i <= '1';
                when 7242 => sda_i <= '1';
                when 7243 => sda_i <= '1';
                when 7244 => sda_i <= '1';
                when 7245 => sda_i <= '1';
                when 7246 => sda_i <= '1';
                when 7247 => sda_i <= '1';
                when 7248 => sda_i <= '1';
                when 7249 => sda_i <= '1';
                when 7250 => sda_i <= '1';
                when 7251 => sda_i <= '1';
                when 7252 => sda_i <= '1';
                when 7253 => sda_i <= '1';
                when 7254 => sda_i <= '1';
                when 7255 => sda_i <= '1';
                when 7256 => sda_i <= '1';
                when 7257 => sda_i <= '1';
                when 7258 => sda_i <= '1';
                when 7259 => sda_i <= '1';
                when 7260 => sda_i <= '1';
                when 7261 => sda_i <= '1';
                when 7262 => sda_i <= '1';
                when 7263 => sda_i <= '1';
                when 7264 => sda_i <= '1';
                when 7265 => sda_i <= '1';
                when 7266 => sda_i <= '1';
                when 7267 => sda_i <= '1';
                when 7268 => sda_i <= '1';
                when 7269 => sda_i <= '1';
                when 7270 => sda_i <= '1';
                when 7271 => sda_i <= '1';
                when 7272 => sda_i <= '1';
                when 7273 => sda_i <= '1';
                when 7274 => sda_i <= '1';
                when 7275 => sda_i <= '1';
                when 7276 => sda_i <= '1';
                when 7277 => sda_i <= '1';
                when 7278 => sda_i <= '1';
                when 7279 => sda_i <= '1';
                when 7280 => sda_i <= '1';
                when 7281 => sda_i <= '1';
                when 7282 => sda_i <= '1';
                when 7283 => sda_i <= '1';
                when 7284 => sda_i <= '1';
                when 7285 => sda_i <= '1';
                when 7286 => sda_i <= '1';
                when 7287 => sda_i <= '1';
                when 7288 => sda_i <= '1';
                when 7289 => sda_i <= '1';
                when 7290 => sda_i <= '1';
                when 7291 => sda_i <= '1';
                when 7292 => sda_i <= '1';
                when 7293 => sda_i <= '1';
                when 7294 => sda_i <= '1';
                when 7295 => sda_i <= '1';
                when 7296 => sda_i <= '1';
                when 7297 => sda_i <= '1';
                when 7298 => sda_i <= '1';
                when 7299 => sda_i <= '1';
                when 7300 => sda_i <= '1';
                when 7301 => sda_i <= '1';
                when 7302 => sda_i <= '1';
                when 7303 => sda_i <= '1';
                when 7304 => sda_i <= '1';
                when 7305 => sda_i <= '1';
                when 7306 => sda_i <= '1';
                when 7307 => sda_i <= '1';
                when 7308 => sda_i <= '1';
                when 7309 => sda_i <= '1';
                when 7310 => sda_i <= '1';
                when 7311 => sda_i <= '1';
                when 7312 => sda_i <= '1';
                when 7313 => sda_i <= '1';
                when 7314 => sda_i <= '1';
                when 7315 => sda_i <= '1';
                when 7316 => sda_i <= '1';
                when 7317 => sda_i <= '1';
                when 7318 => sda_i <= '1';
                when 7319 => sda_i <= '1';
                when 7320 => sda_i <= '1';
                when 7321 => sda_i <= '1';
                when 7322 => sda_i <= '1';
                when 7323 => sda_i <= '1';
                when 7324 => sda_i <= '1';
                when 7325 => sda_i <= '1';
                when 7326 => sda_i <= '1';
                when 7327 => sda_i <= '1';
                when 7328 => sda_i <= '1';
                when 7329 => sda_i <= '1';
                when 7330 => sda_i <= '1';
                when 7331 => sda_i <= '1';
                when 7332 => sda_i <= '1';
                when 7333 => sda_i <= '1';
                when 7334 => sda_i <= '1';
                when 7335 => sda_i <= '1';
                when 7336 => sda_i <= '1';
                when 7337 => sda_i <= '1';
                when 7338 => sda_i <= '1';
                when 7339 => sda_i <= '1';
                when 7340 => sda_i <= '1';
                when 7341 => sda_i <= '1';
                when 7342 => sda_i <= '1';
                when 7343 => sda_i <= '1';
                when 7344 => sda_i <= '1';
                when 7345 => sda_i <= '1';
                when 7346 => sda_i <= '1';
                when 7347 => sda_i <= '1';
                when 7348 => sda_i <= '1';
                when 7349 => sda_i <= '1';
                when 7350 => sda_i <= '1';
                when 7351 => sda_i <= '1';
                when 7352 => sda_i <= '1';
                when 7353 => sda_i <= '1';
                when 7354 => sda_i <= '1';
                when 7355 => sda_i <= '1';
                when 7356 => sda_i <= '1';
                when 7357 => sda_i <= '1';
                when 7358 => sda_i <= '1';
                when 7359 => sda_i <= '1';
                when 7360 => sda_i <= '1';
                when 7361 => sda_i <= '1';
                when 7362 => sda_i <= '1';
                when 7363 => sda_i <= '1';
                when 7364 => sda_i <= '1';
                when 7365 => sda_i <= '1';
                when 7366 => sda_i <= '1';
                when 7367 => sda_i <= '1';
                when 7368 => sda_i <= '1';
                when 7369 => sda_i <= '1';
                when 7370 => sda_i <= '1';
                when 7371 => sda_i <= '1';
                when 7372 => sda_i <= '1';
                when 7373 => sda_i <= '1';
                when 7374 => sda_i <= '1';
                when 7375 => sda_i <= '1';
                when 7376 => sda_i <= '1';
                when 7377 => sda_i <= '1';


                --when 250*1    => sda_i <= '0'; -- START
                --when 250*2    => sda_i <= '1'; -- ADDR[7]
                --when 250*3    => sda_i <= '0'; -- ADDR[6]
                --when 250*4    => sda_i <= '1'; -- ADDR[5]
                --when 250*5    => sda_i <= '0'; -- ADDR[4]
                --when 250*6    => sda_i <= '0'; -- ADDR[3]
                --when 250*7    => sda_i <= '1'; -- ADDR[2]
                --when 250*8    => sda_i <= '1'; -- ADDR[1]
                --when 250*9    => sda_i <= '1'; -- ADDR[0]
                --when 250*10   => sda_i <= '0'; -- ACK
                --when 250*11   => sda_i <= '0'; -- DATA[7]
                --when 250*12   => sda_i <= '0'; -- DATA[6]
                --when 250*13   => sda_i <= '0'; -- DATA[5]
                --when 250*14   => sda_i <= '0'; -- DATA[4]
                --when 250*15   => sda_i <= '0'; -- DATA[3]
                --when 250*16   => sda_i <= '0'; -- DATA[2]
                --when 250*17   => sda_i <= '0'; -- DATA[1]
                --when 250*18   => sda_i <= '0'; -- DATA[0]
                --when 250*19   => sda_i <= '0'; -- ACK
                --when 250*20   => sda_i <= '0'; -- DATA[7]
                --when 250*21   => sda_i <= '0'; -- DATA[6]
                --when 250*22   => sda_i <= '0'; -- DATA[5]
                --when 250*23   => sda_i <= '0'; -- DATA[4]
                --when 250*24   => sda_i <= '0'; -- DATA[3]
                --when 250*25   => sda_i <= '0'; -- DATA[2]
                --when 250*26   => sda_i <= '0'; -- DATA[1]
                --when 250*27   => sda_i <= '1'; -- DATA[0]
                --when 250*28   => sda_i <= '0'; -- ACK
                --when 250*29   => sda_i <= '0'; -- DATA[7]
                --when 250*30   => sda_i <= '0'; -- DATA[6]
                --when 250*31   => sda_i <= '0'; -- DATA[5]
                --when 250*32   => sda_i <= '0'; -- DATA[4]
                --when 250*33   => sda_i <= '0'; -- DATA[3]
                --when 250*34   => sda_i <= '0'; -- DATA[2]
                --when 250*35   => sda_i <= '1'; -- DATA[1]
                --when 250*36   => sda_i <= '0'; -- DATA[0]
                --when 250*37   => sda_i <= '0'; -- ACK
                --when 250*38   => sda_i <= '0'; -- DATA[7]
                --when 250*39   => sda_i <= '0'; -- DATA[6]
                --when 250*40   => sda_i <= '0'; -- DATA[5]
                --when 250*41   => sda_i <= '0'; -- DATA[4]
                --when 250*42   => sda_i <= '0'; -- DATA[3]
                --when 250*43   => sda_i <= '0'; -- DATA[2]
                --when 250*44   => sda_i <= '1'; -- DATA[1]
                --when 250*45   => sda_i <= '1'; -- DATA[0]
                --when 250*46   => sda_i <= '0'; -- ACK
                --when 250*47   => sda_i <= '0'; -- DATA[7]
                --when 250*48   => sda_i <= '0'; -- DATA[6]
                --when 250*49   => sda_i <= '0'; -- DATA[5]
                --when 250*50   => sda_i <= '0'; -- DATA[4]
                --when 250*51   => sda_i <= '0'; -- DATA[3]
                --when 250*52   => sda_i <= '1'; -- DATA[2]
                --when 250*53   => sda_i <= '0'; -- DATA[1]
                --when 250*54   => sda_i <= '0'; -- DATA[0]
                --when 250*55   => sda_i <= '1'; -- NACK
                --when 250*56   => sda_i <= '0'; -- STOP              
                --when 250*57   => sda_i <= '1'; 
                when others => sda_i <= sda_i;
            end case;
        end if;
    end process;



end architecture;